class c_40_1;
    integer i = -5;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_40_1;
    c_40_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00011z01zx01x0zxz01zx1xzx0xz0x0zxzxzxxzzzzxxxxzxxxxzxxzxzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_664_1;
    integer i = 664;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_664_1;
    c_664_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1xzxxx0zz0x11x00001z0z01x0z111zxxzxzxzzxzzxzxzzxxzzxzzxzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1870_1;
    integer i = -310;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1870_1;
    c_1870_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "011zxx10zx01z1010z1xxzz101x11001zxzxzxzzxzzxzxzxzxzzzxxxzxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2063_1;
    integer i = -342;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2063_1;
    c_2063_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx1z00001z1110010xxxzxx0001x10zxzxxzzxzxzzzxxzzxzxxzxzxxzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

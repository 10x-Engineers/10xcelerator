class c_2718_1;
    integer i = -451;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2718_1;
    c_2718_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z00xxzxxxz0x0z01x0zzzzxxxxx0xxzxzxzzzzzzxzzzxxzzzxzxxxxzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3038_1;
    integer i = -505;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3038_1;
    c_3038_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00000101x0xxz0zz0xx001xx0zxxzxxzzxzxzxxxzxzxxxzzxzxzxzxxxxzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_370_1;
    integer i = 370;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_370_1;
    c_370_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zx01zxxxzxz100z0x00x0x0xz0xzz0xxzxzzxzzzxzxxxxzxzzzxxxxzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

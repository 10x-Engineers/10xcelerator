class c_2023_1;
    integer i = -336;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2023_1;
    c_2023_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z10zxz1zzz00x10zzz0xxx0101zz1101xxzxzzxxxxxxxzzzzxxxxxzxxxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

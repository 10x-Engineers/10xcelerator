class c_478_1;
    integer i = 478;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_478_1;
    c_478_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1100xx01001zxx1xxxxz01zz1z00x1zzxxzxzzzxzxzxxxzxzxxxxzxxzxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

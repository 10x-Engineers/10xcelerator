class c_2958_1;
    integer i = -491;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2958_1;
    c_2958_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x11zzx000x0zx0zx0x1xzxx11x1x000zxzxxzzzzxzzzxzzxxxxzzxzzzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_154_1;
    integer i = -24;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_154_1;
    c_154_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zzz0x0z0x00x010z11zxz00z0zx0zxzzzzzxxxxxzxxxxxxxxzzzzzxxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_127_1;
    integer i = -20;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_127_1;
    c_127_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0z1z11zz0x01000x001xzxz0000zzzzzxxxxzxzxxzxzzxzzxxxzxxzzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1717_1;
    integer i = -285;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1717_1;
    c_1717_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00z1xxzxz0zxx0z0z00x1x1zzzxz0x0zzzxzxzzzxxxxxzzzxxxxxxxzxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

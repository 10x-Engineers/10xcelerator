class c_129_1;
    integer i = -127;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_129_1;
    c_129_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxx11xzx0xz011zx1zx0zzzz00z1zx0zxzzxxxzzzxxxxxzxzzzxxzxzzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

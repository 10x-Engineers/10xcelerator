class c_3327_1;
    integer i = -553;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3327_1;
    c_3327_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z0zzz0xx0x1xxz1110xxx100xzx1zxzzxzxzxzzzxzzxxxxxzzxxxzxxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_647_1;
    integer i = -106;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_647_1;
    c_647_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0010x001zz1z110xx01zzx0x000xzzzzxxxxxxzzzzxxxxzxxxzxzzxxzzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1765_1;
    integer i = -293;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1765_1;
    c_1765_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xzxz0x1001xz00z00xzzzxzzz1zzz0xxxzzzxzzxzzxzzxzxzxxxxxzzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2060_1;
    integer i = -342;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2060_1;
    c_2060_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x1xzx1110zz1z01010x000z1100x11zzzzzxxxzxxxzxxzxzxxxzxxzxxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

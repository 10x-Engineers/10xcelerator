class c_2231_1;
    integer i = -370;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2231_1;
    c_2231_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0xzxx00xxx01z0zzxxz0zzz1x0xx0zzxxzxzzzxxxzxxxxxxxzzzxzzxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

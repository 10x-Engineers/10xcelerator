class c_650_1;
    integer i = 650;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_650_1;
    c_650_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xxzx11zzzx0x1z0xx1xz001zzxx1zzxzxzzzzzxxxzzxzxzxxxxzzxzxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2897_1;
    integer i = -481;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2897_1;
    c_2897_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxx1z1zxz0zxx1z000000zzx11101zxxzxzxzzxxxzzxzzzxxxzxzzzzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_716_1;
    integer i = -118;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_716_1;
    c_716_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0100xz1x010x1010zzz0z0001z110010zxxzxxxxxxxxxzzzzxxxxxzzxzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

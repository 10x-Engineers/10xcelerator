class c_2795_1;
    integer i = -464;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2795_1;
    c_2795_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000xzxzx11zxzzzzxz0011xx00z0z0z1xxxxzxxzxxxxzzxxzxzzzzzxxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_775_1;
    integer i = -128;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_775_1;
    c_775_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z1000zzz011000x01001zzxzxxx1xzxxxxxxzzzxzxxzzzzzzzzxzxzzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2107_1;
    integer i = -350;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2107_1;
    c_2107_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010zzz01z00z0xxzz01zz0xz10z10110zxzzzxzzxzxxxzzzxzzzzzzxxzzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

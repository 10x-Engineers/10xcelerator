class c_402_1;
    integer i = 402;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_402_1;
    c_402_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110z0xx10x0x1z0z11x0z1x0xz01x1x1zxxxzxzxxxzxzzxzxzzzxxxxzzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

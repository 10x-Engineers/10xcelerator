class c_644_1;
    integer i = -106;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_644_1;
    c_644_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxx1x00x0xx00xzxz10xx0xzx11z10xxxxxzzzxzxzzzzzxzxxzxxxxxxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_580_1;
    integer i = -578;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_580_1;
    c_580_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110x1xzzxzz1xxz1z01zx11x1xz00101xzzzxxxzxzxxzzxzxzzxzxxzxzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2314_1;
    integer i = -384;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2314_1;
    c_2314_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1110zxzx0xxxz0x01zz0zz0zz10xzxzzzzxxxzzxzzxzzxzxxzzxxzxzzxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

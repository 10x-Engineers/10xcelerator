class c_1225_1;
    integer i = -203;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1225_1;
    c_1225_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xz0110z1zzxzz1zz0x10z1x0z0x1xxzzxxzzxzzzxzxzzzzzzzxxxzzxxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_294_1;
    integer i = -292;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_294_1;
    c_294_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz111x0xx0x1z101xxxx100z0zxxz10xxzzxzxzxxxzxxzxzzxxxzzxxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_688_1;
    integer i = 688;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_688_1;
    c_688_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x11z0zzzz0xx0zz0001x0x11xzxzx0xzzxzxzxxxxzxzzxxzzzzxzzzzzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_934_1;
    integer i = -154;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_934_1;
    c_934_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxx011zxxx0x1zx0xxx0x0x001xxz00zxxxzxxxxxxxxzxzzzzzzxzzzzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

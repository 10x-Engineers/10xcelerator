class c_1381_1;
    integer i = -229;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1381_1;
    c_1381_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1zxxxzxz01zz0z100xzx111010xx1xxzxxzzxzxzzxzzzxxzzzxzxxxzzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1505_1;
    integer i = -249;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1505_1;
    c_1505_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z100zx0z011zxxxxz10x001xzz000xxzxzxxzxxxzzzxxzxzxxxzzxxxzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

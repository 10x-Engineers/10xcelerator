class c_926_1;
    integer i = -153;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_926_1;
    c_926_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1z100xz1xxzzx111zzzx0x1zz1zx0zzxxxxzxxzxxxxzxzzxzzxxzzzzxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_482_1;
    integer i = -79;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_482_1;
    c_482_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz0z010z1x101zz000zzzz11z1101xzzzxzzxzxxzxxxxxzzzzzxxzzzzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2810_1;
    integer i = -467;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2810_1;
    c_2810_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010zz1z111zxz1x1xxxzx0zzxz10z0z0xzzxzxxzxxxxxxxzzxzxxzzzzxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2340_1;
    integer i = -388;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2340_1;
    c_2340_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxzx11x1x000xxzz0x0z1x0xz01x00xxzxzxzxzzzzzxxzxzzzxzzzzzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1762_1;
    integer i = -292;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1762_1;
    c_1762_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x111xz1z1z1z1z0xzz111111xxz1zxzxxxxxzzzzxxzxxzzxzxxxzxxzxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

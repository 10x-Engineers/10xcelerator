class c_796_1;
    integer i = -131;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_796_1;
    c_796_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x0z0xz1111zzx1z1z101z0xx1zxxx1zxzzxzzxzzxxzzxzxzzxzxzzxzxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

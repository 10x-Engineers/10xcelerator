class c_1242_1;
    integer i = -205;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1242_1;
    c_1242_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx101zzx01011z1zz1zz0zzx0x1z00x0xzzzxxxxzzzxxzzxxzzxxxzzzxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_661_1;
    integer i = -659;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_661_1;
    c_661_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z001x1zxzzx1x0z01z0zxzxzxx1z11zxxxzzxzzxxzxxzzxzxzxxzzzxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1971_1;
    integer i = -327;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1971_1;
    c_1971_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z10x1110xxx110zz0zx10110zxzxx1xzxzxzzzxzxzxxxxxzzxzzxzzxxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

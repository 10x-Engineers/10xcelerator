class c_594_1;
    integer i = 594;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_594_1;
    c_594_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxz1zz0xxzxzzx1xz010zz0xx10x01xxzzxxzxxzzxxxxxxzzzzzzxxxzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

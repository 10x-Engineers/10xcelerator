class c_460_1;
    integer i = -458;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_460_1;
    c_460_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxz100110x1x1xzzxz1xzzxzxxzzx10zzzxzxxxxxzxxxzxxzxxzzxxzxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_299_1;
    integer i = 299;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_299_1;
    c_299_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz11xz10zxzx1zxzz1zxzx10xzzx00z1zxzxzxxxxzxzzzxzzxxzxzxzxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

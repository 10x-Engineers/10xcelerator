class c_424_1;
    integer i = -69;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_424_1;
    c_424_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz10x1xzz01x1zzz0xz0z0011z0xx001zzzzzxxzzxxzxxxxzzzzxzzxzzzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2035_1;
    integer i = -338;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2035_1;
    c_2035_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x1z1z1xx01xzxzzx0zx1z1z0zx0z010zxzzzxzxxzxzxzzzzxzzxzzxxzzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_473_1;
    integer i = 473;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_473_1;
    c_473_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01xzz1z01x000x10x11xxz11zzxz0z1zzzzxzxzxzxzzxzxzxzzzzxzxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_130_1;
    integer i = -20;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_130_1;
    c_130_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11101zx1z0zzz01x1xz00xx1011zzzxzzxzxxxzxxxxxxzxzzzzxzzxzzzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_678_1;
    integer i = 678;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_678_1;
    c_678_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xx0z1xxzx0zxxx111xxxz1z1xxz0zxzxxzzzzxxxxxzxxzzzxzxxzzzzxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_690_1;
    integer i = -113;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_690_1;
    c_690_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0xz1011z0x0xxz110111z01xzzx000zxzxzxzxxzxxxzxxxzxzxzzzxxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_321_1;
    integer i = -319;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_321_1;
    c_321_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0101xz10111x001z0z111z0xx00x0x1xxzzxzxxxxxzxxxzzxzxzxzxzxxxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

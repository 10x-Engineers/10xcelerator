class c_113_1;
    integer i = 113;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_113_1;
    c_113_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0x11z1x11z11x00xx011x01z110xxxxzxxzxxxxxxxxxzxxxzzzxxzzxzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

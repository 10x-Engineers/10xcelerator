      `define input_size 16
      `define input_matrix_size 12
      `define output_size 32
      `define bias_size 32
      `define kernel_size 5
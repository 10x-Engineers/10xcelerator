class c_2981_1;
    integer i = -495;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2981_1;
    c_2981_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzzzzz0z0xz1z0x00x1110z1111zz10zxzxxzzzxxzzxzxxxxzzzzxxxxzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2061_1;
    integer i = -342;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2061_1;
    c_2061_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz0zxxz11z00111xx1zzz011100zz00zxzzzzxxzzxzxxxxzzzzxzzxxzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

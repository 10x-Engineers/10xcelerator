class c_418_1;
    integer i = -68;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_418_1;
    c_418_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzx10x111zzz01z1xxxzz0z0z1z01zxxxxzxxxxxxzxzzxzzzxzzxzxxzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

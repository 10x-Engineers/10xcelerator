class c_256_1;
    integer i = -254;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_256_1;
    c_256_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz00z0x00xz01zzzxx01z10x00100xzzxzzzxzzzxxzxzxxzzxxxxzxxzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_754_1;
    integer i = -752;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_754_1;
    c_754_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxx0xzzz000xzx0111z0zz1x01z01xxxzzzzzxzzzzzzxxxxzzxzxxzzzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1014_1;
    integer i = -167;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1014_1;
    c_1014_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzz01x0xz0011x1x0x11xx10zx011zxxxzxzzzzzxxzxxxxxzzxxzxzxzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_699_1;
    integer i = 699;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_699_1;
    c_699_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "100001zzx0z1xz1z0xxzx0xzzzzxxzxxzzzxzzzzzxzxzzxxzzzzzxzzxzzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

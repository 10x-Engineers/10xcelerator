class c_241_1;
    integer i = -239;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_241_1;
    c_241_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zx0010111zxz0001xxx1111zz1zxx11xzxzzxxxxzzxzzzxzxxzxzxxzzxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3360_1;
    integer i = -558;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3360_1;
    c_3360_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zxx01zzx1z00x1zx11z1x11xz0z1zxzzzzxxzxzxzxzzzxzxxxxzxxzxzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

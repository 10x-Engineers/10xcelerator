package include_pkg;

  import uvm_pkg::*;



   

`include "uvm_macros.svh"



`include "Seq_item.sv"
`include "Seqr.sv"
`include "Sequence.sv"

`include "Driver.sv"
`include "Monitor.sv"
`include "Agent.sv"

`include "Environment.sv"
`include "Scoreboard.sv"
`include "Test.sv"

endpackage
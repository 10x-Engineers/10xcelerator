class c_973_1;
    integer i = -161;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_973_1;
    c_973_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzx0xx01x1x0x1x0x0x0111z1zx01xxzxxzxzxzxxxxxxxxxxzzxxxxxxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_578_1;
    integer i = 578;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_578_1;
    c_578_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01x100zzz11z010xxx1xxx0x1x01x1zxxzxzzxxzxzxzzxxzzxzxzxxzzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

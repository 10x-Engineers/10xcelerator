class c_483_1;
    integer i = 483;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_483_1;
    c_483_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z11z1xxzz011xxzz1zz100x0x011zzzzzzxzzxxxxzzzzxzxxzxxzzzzxxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_344_1;
    integer i = -342;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_344_1;
    c_344_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x1zz0z1z0zzx011zz0001001xx1z00zzzzzzzxzzzxxzzzxzxxzxzxxzxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2884_1;
    integer i = -479;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2884_1;
    c_2884_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxzxx00z00x0xxzxzxxzz1001z1x10xzzxzxxzxzxzxzxzxxzxzxxxzxxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

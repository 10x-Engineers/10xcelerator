class c_1487_1;
    integer i = -246;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1487_1;
    c_1487_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0010zzzzx0x00xzzzx1x0zz01x1zxxxxzzzxxxxzxxzxzxxxzxxxzxxzzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_654_1;
    integer i = -107;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_654_1;
    c_654_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzxz10011x0x1zxx1x01zzx0z00x10zzxxxxzxzxxxxxxxxzzxzzzxzxxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

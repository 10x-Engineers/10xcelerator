class c_65_1;
    integer i = -63;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_65_1;
    c_65_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000xzzxxx0xx00zzxxx100zx1xxx1x1zzxxxzxxzxxzxzzzzzzxzzxzxxxxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2359_1;
    integer i = -392;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2359_1;
    c_2359_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101z0xxxz00x1z1x0xxzxz10x101z0z0zxzxzzxzzzxxzxzxxxxzxzxxzzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1603_1;
    integer i = -266;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1603_1;
    c_1603_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz01xxzxxz1zzxx0xz01zxx100zx10xxxzzxxzxzzzzzzxzzxxzzzzxzzxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

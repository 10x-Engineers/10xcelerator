class c_1734_1;
    integer i = -287;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1734_1;
    c_1734_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x101xz000xx100z11zzz100100z1xxxzxzxxzzxxzxzzxxxxzzxxzxxzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

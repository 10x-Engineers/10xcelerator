class c_432_1;
    integer i = -430;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_432_1;
    c_432_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxxzz011zxz11010xzxxzxx1zx1x10zxxxxzzzzzzzzzxxxxzzxzxxzzzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

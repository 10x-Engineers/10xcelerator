class c_2280_1;
    integer i = -378;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2280_1;
    c_2280_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxzx00z01x0xzz0zzz1101xx10111zxxxzzzxzxzxzzxxzxxxzzzzzzzxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2876_1;
    integer i = -478;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2876_1;
    c_2876_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z111zz1xxxxzx1xx1zxxx101zxx1xzxxzzxzxzxxxzzxzxzzxzxzzxxzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_297_1;
    integer i = -48;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_297_1;
    c_297_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xzzzxz001x0z0x1x0xxz01xx0x110xxzxxxzxzzxxxxzxzzzxxzxzzxzzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_250_1;
    integer i = 250;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_250_1;
    c_250_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxx1x1xxzxx1x0xz101z010011z0xx1xxxxzzzzxxzzxxxzzxxxzxxxzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_181_1;
    integer i = 181;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_181_1;
    c_181_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1z1xx0xxz0z01x000z1zxxx101zz0zxxzxxxxxzxzzzxzxxzzzxzxzzzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

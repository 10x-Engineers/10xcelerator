class c_1368_1;
    integer i = -226;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1368_1;
    c_1368_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx1xx0z0110z110x1z0xz1zxzzxzz011zxxzxzzxxxzzxzzxxxxzzzxzxzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_701_1;
    integer i = 701;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_701_1;
    c_701_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z1zxz00111z11111zzz1z1z11z110zxxxzzzzzzzxxzzzzzxxxzxxzxxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3308_1;
    integer i = -550;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3308_1;
    c_3308_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zzzx0z00xx1z1010x0x1z1z1z0z1zzzzzzxzxxxzxxxzxzzzxxxxxxxxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3410_1;
    integer i = -567;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3410_1;
    c_3410_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z01111zx1z10x0zz0x01zzxxz1xzx1xxxxxzxxxxzzxzzxxxzzxzxxzxxxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1963_1;
    integer i = -326;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1963_1;
    c_1963_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x111xzxxzz000011zxx01x001zxxx0z0xxxxxxxzxzxzzxxxzxzzxxxxzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2867_1;
    integer i = -476;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2867_1;
    c_2867_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1xx0z010zz10zxxzxxz1zx1z100xxxzzzxxxzxzxxzzzzzzzzxxxxzzxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

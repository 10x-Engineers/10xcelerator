class c_2638_1;
    integer i = -438;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2638_1;
    c_2638_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z11zzxx001xzx1xxz1x0xxx1z0100zzxzxzxxxxxxzxzxzzzzzxzxzzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

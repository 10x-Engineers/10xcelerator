class c_1192_1;
    integer i = -197;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1192_1;
    c_1192_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzz1x0xxz1xxx0011z1zzx1zxzxz11zzzzxzzzxxzzzxxxzxxzzzzxzxxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_768_1;
    integer i = 768;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_768_1;
    c_768_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z01xzz00z0000zxzzxxz10xx01z1xzzxzzxxzzzxzxzzxxzzzzxxzzxxxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_908_1;
    integer i = -150;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_908_1;
    c_908_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1zzxxxxxz11xxxx11xxx10xxx00zxzzxxzxxzxxxzzzxzxzxzzxzxzxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2520_1;
    integer i = -418;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2520_1;
    c_2520_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01x1x0xxzx0zx1zz001001z000zx0x0zzzzxzxxzzzxxzxxzxzxzzxxzzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

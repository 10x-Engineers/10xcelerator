class c_3084_1;
    integer i = -512;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3084_1;
    c_3084_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x1xx10zzzx1xx0xxxx1z00001zxzx0xzzxxxxxxxzzzzzxzzzxzxzzxzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1513_1;
    integer i = -251;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1513_1;
    c_1513_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1xzz1xzzz01xzz101xx00z1zz11zzzxxxxxzzxxzxxzzzzzzzzzzxzzzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_396_1;
    integer i = -64;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_396_1;
    c_396_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xzx0100x1xz0zzzx00zxzx0z0zxzx11xxxxzxxxzxzzzxxzxxzxxzzxzzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1735_1;
    integer i = -288;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1735_1;
    c_1735_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzxzz11z0zxz1z1110z100xzx0zzz01zxxxxzzxzxxxxxxzzxzzzxxxxzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

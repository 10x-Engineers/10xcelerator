class c_1688_1;
    integer i = -280;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1688_1;
    c_1688_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz110x010xz1000x0zz01100000xz001xxzzxxxzxxxzzzxzxzzxxzxxxxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

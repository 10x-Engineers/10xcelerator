class c_1968_1;
    integer i = -326;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1968_1;
    c_1968_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zz0101101001001100zx1x0z0xzzx0xzzzzzxzzzzzzzzxzxxzzxzxxzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_742_1;
    integer i = -122;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_742_1;
    c_742_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x0xxx010z01xxz1x0x1z0zxxxzzxx0zxzzzzzxxzxzzzxxzxzzzxzxxxxxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

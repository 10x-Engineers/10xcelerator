class c_2928_1;
    integer i = -486;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2928_1;
    c_2928_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xz11z000xxzx1001xzx0zx111zz1xzzxxxzxxzzzxxxxxzzxxxxxxxxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1633_1;
    integer i = -271;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1633_1;
    c_1633_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x100xxxzx1z0z10100zx0000110xz1x0zzxzxzxxzxxzzxzxxxxxzxxxzzxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

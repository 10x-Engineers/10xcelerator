class c_2538_1;
    integer i = -421;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2538_1;
    c_2538_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xx0100xx10zx010z11xzzx1zx0x0xzxzxzxxzzzxzxxxzxzzzzzzzzxzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_847_1;
    integer i = -140;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_847_1;
    c_847_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz1zx1xx0xzzz001xzz1xz0zx1x1xx0zxxzxxxxzxxzzxzxxzxzxzzxxzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_215_1;
    integer i = 215;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_215_1;
    c_215_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x0z00100110zxz1111xx0x0xzzx0xxzzzzxxzxxzzxzxxxzxzxxzxxzxzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3192_1;
    integer i = -530;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3192_1;
    c_3192_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz0zx0xxx1zxzx1z0zzx0x1z0zx1zx1zxzxzzxxzxxzxxxxxxzxxxzzxzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

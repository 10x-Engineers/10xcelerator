class c_1404_1;
    integer i = -232;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1404_1;
    c_1404_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x10z00z01xx1xz10z00x0zzzzz1x101xxxxxxzzxzxxxxzzzxxxxzzxzxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

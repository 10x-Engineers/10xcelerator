class c_2647_1;
    integer i = -440;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2647_1;
    c_2647_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x0x11xzz10zx1x101zz11zz0101x11xxzzxxzxzxxzxzxzzzxxxxzxzxxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1470_1;
    integer i = -243;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1470_1;
    c_1470_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0xxzzzx000z11100x0010zzz1x0xxxzzzzzxzzzxzzxxxzzxzxzzxxzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1805_1;
    integer i = -299;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1805_1;
    c_1805_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zzx0xx0z00xx01z00x011xzx0z0x00xzxzxxxzxxzzxzxxxzzxxxxzxzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

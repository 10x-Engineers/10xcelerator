class c_34_1;
    integer i = 34;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_34_1;
    c_34_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zx1z11010x11xzz0x01000z000010xzzzzzzxzzzzzxzxzxxxxxxzzxxzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_306_1;
    integer i = -304;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_306_1;
    c_306_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z0z1011z01000xxxz10x1z0zxz000zzzzzxxzzxzzxzxxzxzxxxzzzxzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

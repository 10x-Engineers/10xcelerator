class c_740_1;
    integer i = -738;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_740_1;
    c_740_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxx01z11100xx0xxx111zxxz00010xz0xxxxzxzxzzxxxzxzxzxzzzxxxzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1390_1;
    integer i = -230;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1390_1;
    c_1390_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10x01zx10zz0z101z0xz00x1z0x0x1xxxzxzxzxzzxzxzxzzxzxzxxxxzxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

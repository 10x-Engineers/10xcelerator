class c_686_1;
    integer i = -113;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_686_1;
    c_686_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0z111z11x10010z1x1zxz0zz011xxxxxxxxxxxxxxxxxzzzxzzzxxxxzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_118_1;
    integer i = -18;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_118_1;
    c_118_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz0101x01z000xz1x1100x1zz001zz1zxxxxzzxxzzxxxzxzxxxzxzxzxxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2952_1;
    integer i = -490;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2952_1;
    c_2952_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z1zx0z011zx0x01z011z1z1000x0zzzzzzzxzzzxxzxxzzzxzxxxzzzzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

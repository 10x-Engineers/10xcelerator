class c_1659_1;
    integer i = -275;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1659_1;
    c_1659_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z011zzxzzzzz0x1zxx10101zx0xzz1x1zzzxzxxzxzzxxxzzxzxzxzxzzxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_268_1;
    integer i = 268;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_268_1;
    c_268_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz00100x0000xx01xx0xzx0zzzxzx101xzxxxzzzzxxxzxxzxxzzxzzzzxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

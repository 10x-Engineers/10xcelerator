class c_99_1;
    integer i = -97;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_99_1;
    c_99_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz0zx0x100z00x0zz011z1x10x1z11z1zxxxzzzzxzxzzzxzxxzzzzxzxzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2319_1;
    integer i = -385;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2319_1;
    c_2319_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz10z0z0zzz100xz00xxx1xz1001xz0xzxzxzzzxxxxzxxzzzxzzxzzxxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_912_1;
    integer i = -150;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_912_1;
    c_912_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0001x0z1z0xz101x01z1x11zx10x1z1zxxxxxzxxzzxzxxxzzzzxxzxxzzxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1020_1;
    integer i = -168;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1020_1;
    c_1020_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001zz110100zx1z0zzxzxx00xz11z1z0zxxxxzzzzxzxxxzxzzzxxzxxzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_299_1;
    integer i = -297;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_299_1;
    c_299_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zzxz11x00xxz1x110zx11000x10x10zxzxxzzxzxzxzxzzzzzzzzxzxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1618_1;
    integer i = -268;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1618_1;
    c_1618_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110100z1xzx1z0x1z0xz00xzxz101000xxxxxzzzxzzxzzxxxzxzxxzxzzxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram



interface small_if(input bit h_clk);


//int output_bits= 32; // fr time being hardcoding values 
//int input_bits =16;
        wire [32-1:0] output_port1;
        wire [32-1:0] output_port2;
        wire [32-1:0] output_port3;
        wire [32-1:0] output_port4;
        wire [32-1:0] output_port5;
        wire [32-1:0] output_port6;
endinterface: small_if


class c_145_1;
    integer i = -23;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_145_1;
    c_145_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1101zzxzzxzzzxxx0010xxx0z1xz0zxzxzzzxxzxxxxzzzxxxxxzxxzzxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1887_1;
    integer i = -313;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1887_1;
    c_1887_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10zz10xzz1zxz1x1100z110xzzz1101xxzzxzxxxzzzzzxxzzxzxzzzzzxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

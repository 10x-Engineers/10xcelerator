class c_272_1;
    integer i = 272;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_272_1;
    c_272_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z001xx011zx0zzxzxx0xxz0zxz1xz1x1xzzxzzzzxxzzxzxzxzzzzxzzxzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2178_1;
    integer i = -361;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2178_1;
    c_2178_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z0000xz00z01zxzz01xx0xxx01001zxxxzzzzzzzxzxxzzzzxxxxzxxxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

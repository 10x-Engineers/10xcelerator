class c_3328_1;
    integer i = -553;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3328_1;
    c_3328_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11z0zzzz00011z011xx1x01xzxzx0x10zzzzzzxxxxzxxzzzzzzxxxxxzzxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

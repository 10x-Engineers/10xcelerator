class c_2659_1;
    integer i = -442;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2659_1;
    c_2659_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz11001x00zz011x11zz01000xz0xz1zzxxzzzzxxxzxxzzxzxxxzxxxxzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

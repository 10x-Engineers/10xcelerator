class c_1232_1;
    integer i = -204;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1232_1;
    c_1232_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z1z1010zxxz0100xzz0010xz00010xzxxxzxxzxzzxxxxxzzxxzxzzzxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

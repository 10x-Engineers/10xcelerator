class c_1034_1;
    integer i = -171;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1034_1;
    c_1034_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx111xx1zzz00zxzz11z000zx1zzz111zxxzzxxxxxzzzzxxxzxzzxzxxxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

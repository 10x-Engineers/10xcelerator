class c_658_1;
    integer i = -656;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_658_1;
    c_658_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10xzxx0zx10110x0x101x1xxz01z1x11zxxzzzzzxzxzxzxzzzxzxzzzzxzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

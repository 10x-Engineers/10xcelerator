class c_576_1;
    integer i = 576;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_576_1;
    c_576_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1111x1x0100xx0z11zx0z10x111z0z1xxzzzxzzzxxzxxzxzzxzzzzzzzzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

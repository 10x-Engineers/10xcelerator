class c_3173_1;
    integer i = -527;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3173_1;
    c_3173_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx101xzx0xzzzxzx0zxx1xz0zx1z10xxzxzzzzxzxzxxxxzzxzzxxzzxxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2124_1;
    integer i = -352;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2124_1;
    c_2124_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx011110zz0zxx00xz1x0z00xxzxz111zxxzxxxzxxzxzxxxxzxxxzzzzxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

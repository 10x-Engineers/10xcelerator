class c_1904_1;
    integer i = -316;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1904_1;
    c_1904_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1x10z010x011zx011z0xzx1011x100zzxxzxxzzxxxzzxzxxxxzzzxxxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

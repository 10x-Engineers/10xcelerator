class c_2589_1;
    integer i = -430;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2589_1;
    c_2589_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxxxzxxzx00z1001z0x1z11xzzxxx00zxxxxxzxzzzzxxxzzzxzxxzzzxzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_540_1;
    integer i = 540;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_540_1;
    c_540_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xzzx001xxz1x0xzzzxz100011x110xxzxxxzzxzxxxxzxzzxzxzxxxzxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

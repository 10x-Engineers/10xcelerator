class c_644_1;
    integer i = -642;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_644_1;
    c_644_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxz11zz1x1z0zxx1x000z11xzx000xzxxzxzzxxzzxxzzxxzzxxxxzzxxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

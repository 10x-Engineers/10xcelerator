class c_704_1;
    integer i = -702;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_704_1;
    c_704_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00101z1110x00xx1z00110xz10x00110zxxxzxzxzzxxzzzxzxxzzxzxxzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2931_1;
    integer i = -487;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2931_1;
    c_2931_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzzzzx1100x0xz110xx00xz000zz00zxzzxxzzxzzxxzzzxzzzzzxzzzzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

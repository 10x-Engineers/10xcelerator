class c_3116_1;
    integer i = -518;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3116_1;
    c_3116_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x110x1x0z110z0xz11xxzx1z1z10xzxxxzzxzxzzzxzzxxxxzxxzxxxxxzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

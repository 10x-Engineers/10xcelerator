class c_3199_1;
    integer i = -532;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3199_1;
    c_3199_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1xzzz1100xxzzx010zz0z0x0x10xzxzzxxxzzzxzxxxxzzxzxxzzxxzxxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3288_1;
    integer i = -546;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3288_1;
    c_3288_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x001x10000xx100x1000z0000zx0xxxxxzxzzzzzzxzzzzzxzxzzzxzzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

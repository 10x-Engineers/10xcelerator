class c_47_1;
    integer i = -6;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_47_1;
    c_47_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxzzz00xxxzxzzz1xxzxzzz10xz01xz1xzxzxxzxxxxxzzxzzxzxzzxzzzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

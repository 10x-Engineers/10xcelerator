class c_568_1;
    integer i = -566;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_568_1;
    c_568_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx1zxxzzz1zz110110z1x0x0x0xx00z0xzzxxxzzzzzxzzxzxxzxzzxxzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

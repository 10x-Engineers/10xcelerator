class c_2487_1;
    integer i = -413;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2487_1;
    c_2487_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x0x1z1x00z1zz0z0zxz011x0z0z0xzxzxzzxzxzzzxzzxzzzzxxxzzzxxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1082_1;
    integer i = -179;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1082_1;
    c_1082_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x000z001xxzz1xxzxx01x0xx01x0zxzzxxxxzzzxzzxxxxzzzxxzzzzzxzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_246_1;
    integer i = -244;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_246_1;
    c_246_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zx11z01101zxzxzxz01zzxzzxxz0xx1zzxxzzxzzxxzzzxzzxxzzxxzzzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

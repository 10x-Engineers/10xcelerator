 `include "parameters.svh"

interface small_if(input bit h_clk);


//int output_bits= 32; // fr time being hardcoding values 
//int input_bits =16;
        wire [`OUTPUT_SIZE] output_port;
endinterface: small_if


class c_1604_1;
    integer i = -266;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1604_1;
    c_1604_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00101z1z11zxxxxz0zz1zx1zxx0xxzzzxzzzzxxzxxxxzzxxxxzxzzxzzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_776_1;
    integer i = -774;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_776_1;
    c_776_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101zxxzz0x0z01x00100zxzz01zzzzxzxxxxxzxxzzxzxxxzzxxxxzzzzxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

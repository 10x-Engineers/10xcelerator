class c_649_1;
    integer i = -107;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_649_1;
    c_649_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0000z1z1xzxxz01zxzz1z1zxx0zx0zzxzxzxzxxxxzzxzzzzzxxxzzzxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_622_1;
    integer i = 622;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_622_1;
    c_622_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0z1x1z1x11100z01z110xx10z1z010zxzzzxxzzzzxxzxzzzzzzxxzzxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_278_1;
    integer i = -276;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_278_1;
    c_278_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz11x1x1zxzxzz0xzz01xxxx01zx00z1xzzxzxzxzzxxzzzxzzxzxzzxzzxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

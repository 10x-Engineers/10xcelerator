class c_129_1;
    integer i = 129;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_129_1;
    c_129_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz0x1xxzzx10xxx010z1z0xx110z10zzxxxzxzxxzzzzzzzzxzxxxzxxxxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3086_1;
    integer i = -513;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3086_1;
    c_3086_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzzxzz00110x10xx11111zzxz11z11zxxzxxzzzzzzzzzxxxzzxzxxxxxxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

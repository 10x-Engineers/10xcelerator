class c_1466_1;
    integer i = -243;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1466_1;
    c_1466_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx11x1x1xxx01x01xz1xzxx10010xz1zxxzzxxzzxxzzzzxxzxzxxzzxxxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

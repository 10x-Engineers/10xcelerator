class c_411_1;
    integer i = -67;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_411_1;
    c_411_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzx00z1001zx1xzz00x0zxxxxzx0zx1zzzxzzxxzzxzzxxzxzzzxxzzzxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

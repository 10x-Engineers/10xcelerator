class c_2276_1;
    integer i = -378;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2276_1;
    c_2276_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001x00111z00xx0xz0z110101x011000zzzxzxxxxzxxxxzzzxxxzzzxzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3148_1;
    integer i = -523;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3148_1;
    c_3148_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00xzzz101xx0zxz1xx0xxx01z0z0z0xzzxzxxxzxzzxzzzzzxxxzzxxxzzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1855_1;
    integer i = -308;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1855_1;
    c_1855_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz00xxz11z0xzzxz1111zz1xz1101xzzzzzzxzzxzxxxxxzxzxzzxzzzzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

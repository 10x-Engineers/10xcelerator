class c_1939_1;
    integer i = -322;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1939_1;
    c_1939_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x010x1z1z11z101z0zxz11xz11100x1zxxxxzzxzzzxzxxxzxxzxxzzxxzxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

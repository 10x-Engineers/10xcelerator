class c_364_1;
    integer i = -362;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_364_1;
    c_364_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx1101000xzxz0z1z0zz1xz000zz01xxzxzzzxxzzxxxxxxxzzxzxxxxzzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

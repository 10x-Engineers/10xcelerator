class c_488_1;
    integer i = -80;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_488_1;
    c_488_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzz001xxzz10zxzx00xzxxx1zzx00xz0xxzzxzzzxzzzxzxxxzzzzzzxxzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

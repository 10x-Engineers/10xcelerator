class c_102_1;
    integer i = -100;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_102_1;
    c_102_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "011xxx0x0xz0zz101xx0x100x1xzxzxzxxzxxzzxxxxzzxzxzxzzxxzzxxxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

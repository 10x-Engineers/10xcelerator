class c_464_1;
    integer i = -462;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_464_1;
    c_464_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xz0zz0x1z011011z1010z0x001xzz1xxzzzxzzzzzxxzxzzzxzxzzxxxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

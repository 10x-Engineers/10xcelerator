class c_1502_1;
    integer i = -249;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1502_1;
    c_1502_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001zxzz01zz01x11z01xxx10xz0xzzzzxxzxzzxzzxxxzzzxxzxxxzzxzxzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

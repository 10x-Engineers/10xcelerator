class c_3200_1;
    integer i = -532;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3200_1;
    c_3200_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz1zz1zx1z00zzxz100010z0xxzxx00xzxxxxxzzzxzzxxzzxxxxzxxzzzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1078_1;
    integer i = -178;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1078_1;
    c_1078_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xz0z001xz10zzxx01z11z00z01000zzxzzxxzxzxxzzzxzzzxzzxzxzzxzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

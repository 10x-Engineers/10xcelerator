class c_1388_1;
    integer i = -230;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1388_1;
    c_1388_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x00110x101110001x1110x1zz01z110xxzxzxzzzxzxzxzxzxzzxzzzzxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_460_1;
    integer i = -75;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_460_1;
    c_460_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzzzxx00x1000zxzxz10x0x0x11z01zxzzzzxxxzxxxzzxxzxxzxzzxzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1634_1;
    integer i = -271;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1634_1;
    c_1634_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0000z1x0zz111x101zzx0x1zz0z00000xxxxzzzxxzzzzzzzxzxxzzxxzxzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2008_1;
    integer i = -333;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2008_1;
    c_2008_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz00z01z1x111zzz001xxx1zx00zz00xzzxxzzzzzxzxxxzzzzzxxxxxxxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2102_1;
    integer i = -349;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2102_1;
    c_2102_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xz111zx1x0xz11x011z0xzxzx1110xzxxzxzxzxzzzzzxxxzxxxzzzzxzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2979_1;
    integer i = -495;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2979_1;
    c_2979_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11z1xz10xzxzz0zzzz0101xx110zzxzzzxxzxxxzxxzzxzzxzzxzxxxxzzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_646_1;
    integer i = -644;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_646_1;
    c_646_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xzx10z10z1z1101z0x11x10x0zz0xzxxxxxxzzzzxzzzzxzxzxzxzzzzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

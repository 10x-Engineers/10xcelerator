class c_898_1;
    integer i = -148;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_898_1;
    c_898_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x0zz0zxxzx00x11xz0xzzx1x0zxzx1xxzxzzxzzzzzxzxzzxxxxxxzxzzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1879_1;
    integer i = -312;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1879_1;
    c_1879_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x000010xzz1110zx100xxz011zx01x0xxxzxzzxxzxxzzzzxxxzzzxxxxxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_476_1;
    integer i = 476;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_476_1;
    c_476_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz0100x0x1x01zxx0xz1zxzx0xx11xxxxxzzzxzzzzzxzxzxzxxxzxzxxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

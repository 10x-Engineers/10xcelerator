class c_281_1;
    integer i = -279;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_281_1;
    c_281_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z010xxz00z01z1xxx011000z1xx0xxxxzxxxxzzxxzzzxxzxxxzzxxxxxxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

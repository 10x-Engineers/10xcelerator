class c_1313_1;
    integer i = -217;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1313_1;
    c_1313_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x1xzxz100xz010xzx1xzx0z11z0z11zzzxxxzzxxzzzxzxzzzzxzzzxzzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3270_1;
    integer i = -543;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3270_1;
    c_3270_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0z1z0011xx1zz0xxx0x0x0x01z1zzxzzzzxxzxzzxzzxzxxzzzxxxzzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

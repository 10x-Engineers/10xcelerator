class c_2517_1;
    integer i = -418;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2517_1;
    c_2517_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x000x0xxx1x000zzzxzx1x1110x01x0xzzzzzzzzzxxzzzzzzzxzzzzzxxzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2812_1;
    integer i = -467;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2812_1;
    c_2812_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0000xx00zxx0x00x11x1zx011z0xzzzzxxxzxzzxzxzxxzxxxzzzxzzxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

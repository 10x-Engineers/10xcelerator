class c_773_1;
    integer i = -771;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_773_1;
    c_773_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000z0100x0x1011z00x1z0xz0zxzzxzzzxzzxxzzzzxzzxxxxxxxxzxxzxzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

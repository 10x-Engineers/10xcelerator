class c_2147_1;
    integer i = -356;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2147_1;
    c_2147_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z11zxxzz01x0xz0z10x11z1x11xzx0x1zxzxxxxzzxzxzzzzzxzzzzzxzzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

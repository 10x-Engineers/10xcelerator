class c_66_1;
    integer i = -9;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_66_1;
    c_66_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxzzx10xzz1xzxz0001z0z00xx101zz1zxzxxxxzzzzzxzzxzzzxxzxzzxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_531_1;
    integer i = -529;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_531_1;
    c_531_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z110110xx1zx00zx10z000x011xzx0x1xzxzxxzzxxxzxzxxxzzxxxzxxzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

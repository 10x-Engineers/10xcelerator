class c_385_1;
    integer i = -63;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_385_1;
    c_385_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz101x100001x1xz0zxzxx11zzx1zx0zzxzzzxzzxxxzzxxxzxzzzxzxxxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_619_1;
    integer i = -617;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_619_1;
    c_619_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0x1zxzzz0xz01zzz1zx1x1xx010zxxxxxzxzzzxzxxxxxxxxxxzzxxxzxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

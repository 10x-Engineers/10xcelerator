class c_164_1;
    integer i = -162;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_164_1;
    c_164_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z10zzxxxz10111xxx011zz001z010x1zzzxxzzxzzxxzxxzxxzxxxxxxzxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

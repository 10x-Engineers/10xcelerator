class c_333_1;
    integer i = 333;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_333_1;
    c_333_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x00xzx00zxxzxz1xx11xzz0z1zzxx0xxzxzzxxzzxzzzxzxxzxxxxzzxzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_661_1;
    integer i = 661;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_661_1;
    c_661_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111x00z0x1z0xx11xzxxxxz0xz00x1x0zxzzxxzzxzzzxxxzxxzxxxxzxxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1556_1;
    integer i = -258;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1556_1;
    c_1556_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xz10010xzx110001z1zz101x0zzxx00xzzzxzzzxxzxxzzxzzxxzxzzzxzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_286_1;
    integer i = -46;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_286_1;
    c_286_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxx100z0zzzxxx00z0zx1xz10xx11zzzzxxzxxxxxxxzxzzxxxxxzxxxxxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

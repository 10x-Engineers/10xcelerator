class c_2079_1;
    integer i = -345;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2079_1;
    c_2079_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz1xz00x10xxxz01010xxxx111x1xx0zxzzxzxzzzxxxzxzxxzzzzzxzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_51_1;
    integer i = -49;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_51_1;
    c_51_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0z01zxz0z0zx1x001101z0z1xxzx1zzxzzxzzxzxzxxzzxzzzzzxzzxxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2567_1;
    integer i = -426;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2567_1;
    c_2567_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z100z00zzz1100x000z1xx00xxzzx1zxzxzzxxzxzzxzzzxzzzzxzzzzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

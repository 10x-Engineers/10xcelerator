class c_376_1;
    integer i = 376;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_376_1;
    c_376_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxx00x00x111zzx1xxzzxz0xx01xx00zzxzxzzxzzzxzzzzzxxxxzxzzxxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

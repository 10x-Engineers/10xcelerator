class c_2569_1;
    integer i = -427;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2569_1;
    c_2569_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zz01zzx1xxxxx1110z0z01xz01zzx0zzzzxxzzxxzzxxzxzxxzzzxxxzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3414_1;
    integer i = -567;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3414_1;
    c_3414_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10x0z10zz01z01x0z1xz1zxx000xxzzzxxxxxzzxzxzxzzxxxzxxzxzxzxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

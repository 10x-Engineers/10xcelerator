class c_2657_1;
    integer i = -441;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2657_1;
    c_2657_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzzzzxz11x1010xx110zz00xx0z10zxxzxxzxxzzxxzzzxxzxxzzzzzxzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

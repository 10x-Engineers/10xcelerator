class c_558_1;
    integer i = 558;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_558_1;
    c_558_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "100001x0zx0xxx1xxxxzx0x11x01z0x0zzzxxzzxxzzzzzzxzxxzxxzzzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

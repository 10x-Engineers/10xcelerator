class c_1492_1;
    integer i = -247;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1492_1;
    c_1492_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz00x0zz011z101000zz11xz0zzx10xxxxzzzzzxxzxxzxxxzzzzxxzxxxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_187_1;
    integer i = 187;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_187_1;
    c_187_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1001xx10zz0x10zx0xzx10000xxxzxxxxzzxzzxzxzxzxxxzxzzxxxxxxzzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2175_1;
    integer i = -361;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2175_1;
    c_2175_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzx0001z00xz0zzx1x0zz101z1zz10xzzzzzxzzxzxxxxxzxzxzxzzzzzxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2494_1;
    integer i = -414;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2494_1;
    c_2494_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z1x10z011xzzzz10xx1000z10zx1zzzzzxzxzzzzzxzxxzxxxxzzxxzzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

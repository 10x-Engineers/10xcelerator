class c_2552_1;
    integer i = -424;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2552_1;
    c_2552_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xzx0zx1101000zzz11z010zz1x000zzzzxxzzzzxzxzxxzzxzzzxzxzxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

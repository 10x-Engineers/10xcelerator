class c_492_1;
    integer i = -80;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_492_1;
    c_492_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zz1xx1x00zz00zx010z1z11zzx1x11xzxzzzxxzzzzzxzxzzzxxzxzzxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

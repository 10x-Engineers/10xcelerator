class c_2685_1;
    integer i = -446;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2685_1;
    c_2685_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11z11001zz00x10x001z1z001zx0100xzxxzzxzzzxzzzxzzzzxzxxxxxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_753_1;
    integer i = -751;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_753_1;
    c_753_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz0zxx0z001z00100z1zxzzz11xzx10zzxxxzxzzzzxxzzxxzzzxzzxzxxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

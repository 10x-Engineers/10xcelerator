class c_2782_1;
    integer i = -462;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2782_1;
    c_2782_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x001zx0x1xz1xxx1x101x11zzx1x01xxzzzxzxxxxxxzxzzzzxzzxxxxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_319_1;
    integer i = -317;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_319_1;
    c_319_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010zx1zzx00z0xx1x0x010z10xz11111zzxxzzzxxzzxzzxzzxzzzzzzxxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1948_1;
    integer i = -323;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1948_1;
    c_1948_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x1x001x1zz10011zzz011101z1xzz0xzzxxxzxxzxxxzxzzxxzxxzxxxxxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

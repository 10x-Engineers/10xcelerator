class c_809_1;
    integer i = -133;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_809_1;
    c_809_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzx1xz0xz1x0x110x0x01z0z11z00zxzzxzzxzzxzzzxzxxzzzzxxxzxzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2976_1;
    integer i = -494;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2976_1;
    c_2976_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0xzz000111z111z0zzzx00x100z101zzzxxxxzxxzzzxzzzxzxxzxxxxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_501_1;
    integer i = 501;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_501_1;
    c_501_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z00x001xzx00xz1x00110xzx10xxz1zzxzzzzxzxzxxxxxzxxzzxzzzxxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

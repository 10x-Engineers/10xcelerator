class c_769_1;
    integer i = -127;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_769_1;
    c_769_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z11zz001100zz101xx0x10000x1z10xzzxzzxxxxzzzxzxzzzzzxxzzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

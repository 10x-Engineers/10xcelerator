class c_1817_1;
    integer i = -301;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1817_1;
    c_1817_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz0x1z101z01111xxxxx10x00x111xxxxxxzzzzxzzxxzzxxzzzxzxzzxxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

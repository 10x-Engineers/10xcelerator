class c_1803_1;
    integer i = -299;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1803_1;
    c_1803_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx1z000x1z1x1x001xx1010zx0z00xxzxxzxzzzzzxzxzzzxzxxxxxxxxzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_325_1;
    integer i = -323;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_325_1;
    c_325_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0z11z010x1111101zz1xzx0xzxzz1zzzzxxxzzzxxxzxzzxxzzxzxzzzxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

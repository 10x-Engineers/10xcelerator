class c_2721_1;
    integer i = -452;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2721_1;
    c_2721_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxzz00z1zz0001xz1zzzxx1001zz11zzxxxxxxxzxzxxzxzzzxzzxxzzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_570_1;
    integer i = -93;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_570_1;
    c_570_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "011xz0xxx1z111z10xzzx0z1x01zzzxxzzzxzxxzzxzzxxzxzzzxzzxxxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

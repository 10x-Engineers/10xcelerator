class c_1066_1;
    integer i = -176;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1066_1;
    c_1066_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzxxxzz1001z0x1z101zz01xzx110xzzzxxxzzxxzzzzxxzzzzxzxxxzxxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

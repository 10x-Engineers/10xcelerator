class c_1479_1;
    integer i = -245;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1479_1;
    c_1479_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xxx11011xx1111x1xxxzx1000xz1zxxxxxzzxzxzzxzzzxzzzxzzzzxxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

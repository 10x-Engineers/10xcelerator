class c_717_1;
    integer i = -118;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_717_1;
    c_717_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z01zx10x1z000xzzx0zxz10zzz1z011xzzxxxxxzzzzzzxxzzxxzxzzzzzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_579_1;
    integer i = -95;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_579_1;
    c_579_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzxxzzz1zx0xxz0x00x0x01xzz111xzzxzzzzxzxxxxxxzxxzzzzxzzxxzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

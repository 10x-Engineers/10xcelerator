class c_1677_1;
    integer i = -278;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1677_1;
    c_1677_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zx00xxxz00zxxzzxzz0z0z0x10xzz0zxxzxzxxzxzzzzzzzxzzxzxzzxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3059_1;
    integer i = -508;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3059_1;
    c_3059_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxx00zxz00010000z0z01xx01x010xzzxzxxzzxzxzzxxxzzxzxzxxzxxzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

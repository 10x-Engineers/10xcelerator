class c_1916_1;
    integer i = -318;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1916_1;
    c_1916_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x11zzx00zxzzz011zxzxzz100zzxx1xzxzxzxzzxzxxxzzzxxzxxzxxzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2674_1;
    integer i = -444;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2674_1;
    c_2674_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111z00zx0xxx1111x0xx00z10zz0x1x1zzzxxzxzxxzzzzxxxzzxxzzzxxzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_325_1;
    integer i = -53;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_325_1;
    c_325_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z111001zx0xxxzz1101x101xzxz11x0zzxxxxxxzxzzzzxxzzzxzxzzzxzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_444_1;
    integer i = -442;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_444_1;
    c_444_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzz1x11xz0x11zx01xxzxxx011x00xzzzxxzzxxxxzzxzzzzzxxxzxxxxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

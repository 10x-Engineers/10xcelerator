class c_512_1;
    integer i = 512;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_512_1;
    c_512_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0x11zx1z110z0x1x0011000z1z0xzxzxzxzxzzzxxxzxxzxzxzzzxxzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

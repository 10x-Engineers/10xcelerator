class c_493_1;
    integer i = 493;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_493_1;
    c_493_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzz11010x0zzxz011zzzz1xxxxxz01zzzxzxxzzxxzzzzxzxzxxzxxxxxzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_391_1;
    integer i = -64;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_391_1;
    c_391_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0001x100zzz1x110zzz000x10xz010xzxzxzzxxzzzzxzzzzzzzxxxzxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_581_1;
    integer i = -95;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_581_1;
    c_581_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110x1zxx010x11z11x10xz11z1x00001xxxzzxzxzxzzzzzxzzxzzzzxxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

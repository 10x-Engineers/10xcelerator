class c_379_1;
    integer i = -62;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_379_1;
    c_379_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xx0x1z1z1011zzz0x1x00x0x000z11xzxxxxzxxzxzzzzzxxxxzzxzzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1811_1;
    integer i = -300;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1811_1;
    c_1811_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xz0x110x10x01x01xx0011xxxx0z00zzzzxzzxzzxxzxzzxxzzxxzxxzxzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1098_1;
    integer i = -181;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1098_1;
    c_1098_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110zz1z00zz11zzzxzxzx00101z00100zxxxxxxxxzxzxxzzzzzxzzzzzzxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

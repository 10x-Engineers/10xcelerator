class c_1673_1;
    integer i = -277;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1673_1;
    c_1673_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x1z0x1010zx0x1z0z1x1x1z10xxzz0zzzxzzzzxxxxxxxxzzzzzxxzzzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1508_1;
    integer i = -250;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1508_1;
    c_1508_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zxxz1xz0000xxz1z0xxxxzzz10110zzzxxxzxzxxxzzxxzxxxxxzzzxxzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

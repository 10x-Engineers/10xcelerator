class c_1955_1;
    integer i = -324;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1955_1;
    c_1955_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00xx01x11z11x00zx11111x1x11xxxz0zxzzxzxxxzzzzzxxxxxzxxzxxzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1706_1;
    integer i = -283;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1706_1;
    c_1706_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1xx0xzzxzz1x000z000xx1x11x1xzzxxxxzzxxzxxxzxzxzxzxxzxzzxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

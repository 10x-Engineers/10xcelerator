class c_171_1;
    integer i = -169;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_171_1;
    c_171_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10zxzzzx1zz1xxz1z1x1x0z1z001x0xzzzxzzzxzxzzxxzzzxxzxxzxxxxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_486_1;
    integer i = -79;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_486_1;
    c_486_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0101xzxx0x1z1x10x0zz1xx10x0xxxxzzzzzzxxxzzxzzxzzxxzzzxxzzzxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

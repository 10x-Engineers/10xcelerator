class c_1345_1;
    integer i = -223;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1345_1;
    c_1345_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1xx0zzxzzxxxx1zx0zz0x0xxxx01z1zzzxxxxxxzzxxxzxxxxxxxzzxzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2210_1;
    integer i = -367;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2210_1;
    c_2210_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z0010xxz1xz1x001z1100zzx011x11zxzxxxzxxzzzzzxxxzxxxzzzxzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2077_1;
    integer i = -345;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2077_1;
    c_2077_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z1zxxx001xxz00z1zz11010z10zxz1xxxxzxxxxxxxzxxxxxxxzzxzzxzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1326_1;
    integer i = -219;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1326_1;
    c_1326_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzzx0x1xx1xx000z0xxz0zxz0111zx1zzxxxxxxzxzzxzxxzxxxzxzzxxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

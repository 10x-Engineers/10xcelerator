class c_3111_1;
    integer i = -517;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3111_1;
    c_3111_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00zz1zxz0zz0x1xzxz000zxz01z0100zzzxzzzzxzxxzxxxzxzxxzxxzzzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1907_1;
    integer i = -316;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1907_1;
    c_1907_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xx00xzx01xx00110zzxxx0zxz1010xzzxzxxzzxxzxxzzzxzxzzzzxxzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_155_1;
    integer i = -153;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_155_1;
    c_155_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1x10001zzxxx000000zxx10z100xxx0zzzxxzxxxzxxzzxzxzzzxxxxzzzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

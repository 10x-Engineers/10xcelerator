class c_494_1;
    integer i = -81;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_494_1;
    c_494_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z001zx0001zz11111x0zxx1010110xxxxxzzxxxxzxxxzzzzzxzxxzzxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

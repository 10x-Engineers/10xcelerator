class c_1684_1;
    integer i = -279;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1684_1;
    c_1684_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1100zz1000xz1zx11xx11zx1zxzzzxzzxzzzzzzxzzxzzzzzxzzzzzzzzzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_839_1;
    integer i = -138;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_839_1;
    c_839_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zz0x10z0xz1x11xzx0zzx1z0zxz1xzzzzzzxxzzxzzzxzxxxxxxzxzxzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2857_1;
    integer i = -475;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2857_1;
    c_2857_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z1101xxzxz10x0zxxx1110xzz1101zzxxxzxxzzzxzxxzxzzxzzxxxxxxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

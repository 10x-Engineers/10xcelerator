class c_202_1;
    integer i = 202;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_202_1;
    c_202_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx10xzxxxxzxz10110x0z010z1xz10xxxzxxxxxzxxxxxzzxxxzxxzzzxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_980_1;
    integer i = -162;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_980_1;
    c_980_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzxxz010zxz101x00z001z0zxxxx11zxzzxzxxxxzzxzzxxxzxzzxzxxxzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

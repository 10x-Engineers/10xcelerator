class c_2454_1;
    integer i = -407;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2454_1;
    c_2454_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x00xx0z00zx1z110zzzzz010001z110zxzxzxzzzxxzxxzzzxxzxxzzzzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2332_1;
    integer i = -387;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2332_1;
    c_2332_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01zxx0zx1x1zx000x0zx1zzz10xzzzz1xzzzxzzxxxxxxzzzzxzzxzzzxxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

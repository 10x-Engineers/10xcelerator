class c_2543_1;
    integer i = -422;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2543_1;
    c_2543_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz00zzzz1zzx1zx0x0x0000000100xzzzxxxxxxzzxzxzzzxxzxzxzzzxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

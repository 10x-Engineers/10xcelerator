class c_1738_1;
    integer i = -288;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1738_1;
    c_1738_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "100z001x0zzz11z1010z01zz0x01z0x0zzzzzzzzxxxxzzzzxzzzzzzzxzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

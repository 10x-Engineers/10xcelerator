class c_684_1;
    integer i = 684;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_684_1;
    c_684_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x1xzzz00xz0x10zzz111x1xz0xzxz1xxxzxxxzxxxxzzzxxzxxxxxxxxzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_582_1;
    integer i = -95;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_582_1;
    c_582_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010x10zzzzx01zz1xx1xzx0x01zz1x0zzxzxxxxzxxxzzzxxxzxxxzxzxxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

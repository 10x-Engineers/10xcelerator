class c_716_1;
    integer i = -714;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_716_1;
    c_716_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz01xx0x00x011xz11z0x00100xzz10zzxzzzzzzzxxzxxxxxzzxxxxxxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

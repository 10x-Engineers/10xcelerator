class c_2420_1;
    integer i = -402;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2420_1;
    c_2420_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z11zzxz0z1xzz0zx01xz0zz01z0z01xzxxzzzzzzzzzxzzzxxxzxxxxzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1352_1;
    integer i = -224;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1352_1;
    c_1352_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zxxz101011x111111x0xxzxxz1z0xxzxzxxxzzxxzxxxxzxxxzzzxzzzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

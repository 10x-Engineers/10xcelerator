class c_351_1;
    integer i = -349;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_351_1;
    c_351_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz10001xz00zx1xzxzzzx110x011xx0xzzzzzzxxzzxzzzzzxxxzxzxxzxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

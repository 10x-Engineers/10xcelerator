class c_764_1;
    integer i = 764;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_764_1;
    c_764_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "011x01x011xzz11zzx10x1000xxx1z0zxzxxxxxxzzzzzzzxxzzxxxxzzzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

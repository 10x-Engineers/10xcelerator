class c_1130_1;
    integer i = -187;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1130_1;
    c_1130_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxzx1zz1111xx01011x01xx1xzz11xxzzzzxzzzzxzxxzzzzxxzzxxzzxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

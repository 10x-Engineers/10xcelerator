class c_1244_1;
    integer i = -206;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1244_1;
    c_1244_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx110xz11z00zxxzz1xxx0x1zxx0xz1xxzxxzzzxzxzxxzxzzxzzxxxxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_535_1;
    integer i = -533;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_535_1;
    c_535_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1z110z101zz1z10001xzzzx001x101zxxxzxxzzxzxxzzxzxxzzzzxzxxzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1297_1;
    integer i = -215;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1297_1;
    c_1297_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01z1zz0zx010xxxxz100101zzz1zzzzzxzzzxzxxzxzxxzzxzxxxxzxxzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

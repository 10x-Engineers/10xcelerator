class c_26_1;
    integer i = 26;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_26_1;
    c_26_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0010zx1xxz0zx1zz0xx0xzzx0z01z0xxzxxxxxzzzxzxxxxxzxzxxxxxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

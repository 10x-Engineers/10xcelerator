class c_218_1;
    integer i = -35;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_218_1;
    c_218_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xz1z00xxz0zz0x11110zx1x110011zzxxxxzzxxxxzzzxxxzxxzzxxzzzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1229_1;
    integer i = -203;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1229_1;
    c_1229_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10zx00zzxz1x0xxx00xxzz0xzxz1001xzxzzzxzzzxxxxzzzzxzzxzxxxxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3041_1;
    integer i = -505;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3041_1;
    c_3041_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zxx000zz10x11z0x1xz11z0x1z100zxxxxxxzxxzzxxzzxxzzxxzxxzzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2941_1;
    integer i = -489;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2941_1;
    c_2941_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xx0xzzz000x1000xx0xx010z100z11xxzxzzzzxzxzxzzzxxzxxxzxxzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

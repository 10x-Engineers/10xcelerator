class c_1987_1;
    integer i = -330;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1987_1;
    c_1987_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00x11z00z00x1xz1z1x101zxzzzx0z0zzxxxxzzxxxzxzxzzxxxxxxxxzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3004_1;
    integer i = -499;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3004_1;
    c_3004_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx011zzxzxz1xxz0xzxxxzxz1zxx10x0zzzxxxxxzzxxzzxxxzxzzzzzzzxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_592_1;
    integer i = 592;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_592_1;
    c_592_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1111z1100xxxxzxx0110x1100zx110zzzxzzxxxxzzxzxxxxzzxxxzzxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2733_1;
    integer i = -454;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2733_1;
    c_2733_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0x000xz11z0x1x0111010z01x001z1zzzxzxxxxxxzxzzzxzzzxzzxxzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1742_1;
    integer i = -289;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1742_1;
    c_1742_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01z0xzxz0xzx10xxz0zzz1xxz10zxxzxxxzxzxxzzzzxxxzxzxxxzzxzxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2497_1;
    integer i = -415;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2497_1;
    c_2497_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z11z1zxxxz1zxx001xxx11xz1z010xzzxzzxzzzzxzzxxxxzxxzxxzxzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_344_1;
    integer i = 344;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_344_1;
    c_344_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001zzx1x1100z1100xxxxz11x0z1z0z0xxzxzxzzzxzxzzzxzzzxxxxzzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

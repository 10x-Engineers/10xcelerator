class c_40_1;
    integer i = -38;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_40_1;
    c_40_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zz0x1x01xzx00x01000x1x010xz1xzzzxzxzxxzxzxxzxzxzxxxxxxzzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2240_1;
    integer i = -372;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2240_1;
    c_2240_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xzx101x001z01z1x00zz001z1xz0zzxxzzzzxxxxxxzxzzxzxxxxxzxzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_571_1;
    integer i = -569;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_571_1;
    c_571_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000xxzz11x00xx0xxx0zx01x0xz0x0z0xxxxzzxxxxzzxxzxxxzzxzzzxzzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1202_1;
    integer i = -199;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1202_1;
    c_1202_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z10zzz11111xxz11xxxxz0x11xz1xxxzzxzxzzxxzxxzzxzzxxxzxxzxxzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2523_1;
    integer i = -419;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2523_1;
    c_2523_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1xz000000011111x0110x111z1z001zxzzxzzzzzzzxxzxxzxzxxxzxzzzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1256_1;
    integer i = -208;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1256_1;
    c_1256_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx0zzzz1100x1z10z110x0x011001xzxxxzxxxxzxxzzxzzxzzzxxzzzzxzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1984_1;
    integer i = -329;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1984_1;
    c_1984_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xz01z11x011x10101zxxx0zxxz111xzxzxxzzzzzxzxxxxxxxzxzxxxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

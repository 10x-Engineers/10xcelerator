class c_2729_1;
    integer i = -453;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2729_1;
    c_2729_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1z00x001zz1xxzxz1zx100zzz0x111xxzzzxxxxzzxxxzzzxzxxxxzxzzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

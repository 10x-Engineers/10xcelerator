class c_2934_1;
    integer i = -487;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2934_1;
    c_2934_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x0zx0zz00zxxz100z0x0101xx0111xzzzzxxzxxxzzxxzzzzxxxzzzzzxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

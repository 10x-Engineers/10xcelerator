class c_855_1;
    integer i = -141;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_855_1;
    c_855_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00xzz1001zxz1zzx1xzxx1000x00x0xxxzxxzzzxzzxzzzxzzxxzzxzzzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3345_1;
    integer i = -556;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3345_1;
    c_3345_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzz1011z01xzz1zz0zxz0zz0z11xz11xzzxzxzzxzzzzzzxxxxzzxzxxzzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_383_1;
    integer i = -62;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_383_1;
    c_383_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0xxxzxxxz1zzxx00110x001x0z0xzxzzzxxzxzzzxxxzxxzzxzzxxxxxxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

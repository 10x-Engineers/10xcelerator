class c_641_1;
    integer i = -639;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_641_1;
    c_641_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxxxx0zzzz01x10z0xz0zz01x1x1zz0xxzxxxxzzxxxzzzxxxzzzzzzxzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1264_1;
    integer i = -209;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1264_1;
    c_1264_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01zxxxzz100xzx10z0xx0101zz10z0zzzzzzzxzzxxzxxzxzxxzzzzzxzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3348_1;
    integer i = -556;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3348_1;
    c_3348_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1xx10010x1x0xxxx0110zx00zz1zxzzzzzxxxxxzxxxzxzxzxxxzzzxxzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

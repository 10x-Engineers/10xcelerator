class c_110_1;
    integer i = -17;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_110_1;
    c_110_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz0xz0zzx101x111zz0z000xzx101xzzxzxxxzxxzzzxxxzzxxzxzxzxzzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

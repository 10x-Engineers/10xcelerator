class c_2916_1;
    integer i = -484;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2916_1;
    c_2916_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzxz01x01x01zzx1z100zz100x1zx11xzzxzzzzzxxxxzxzzxzzxzzxxxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_451_1;
    integer i = 451;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_451_1;
    c_451_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xz00zxx001z0001zx11x0zx1xx0x00xzxxxzzzxzxxzzxzzzxxxxzxxzzxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

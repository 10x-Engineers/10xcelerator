class c_1883_1;
    integer i = -312;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1883_1;
    c_1883_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxxzxz011z0zxxzzx0xzx1z1xxx1xz0zzxxxzxzzzzxxxzxxxxxxxzxzzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

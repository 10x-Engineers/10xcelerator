class c_1554_1;
    integer i = -257;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1554_1;
    c_1554_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxzz000100zx111x1zz0100x010x11xxzzzzzzxxzzxxxzzxzzxxxzzxxzxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1281_1;
    integer i = -212;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1281_1;
    c_1281_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xx0xzxz01x10z1xxxxzz0z1zxz011xzxxxzxxzzxzzzzzzxzzxzxxxxxzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3447_1;
    integer i = -573;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3447_1;
    c_3447_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0zx001zz0xzz001zxzx0x1z000xz0xxzzzxzzzxzzxzxzxzxzxzxzzxxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1858_1;
    integer i = -308;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1858_1;
    c_1858_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zxz1xzz0z10xxzxz000xxzzz1xz0xxxzzxxzzzzxzxzxxzxxzxzxxzzzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

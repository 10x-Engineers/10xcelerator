class c_2914_1;
    integer i = -484;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2914_1;
    c_2914_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zxx0xzzz1zx10x1z0zz010xzzz0z01xzzxxzzzxzxxzxzzxxxxzxxxzzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_783_1;
    integer i = 783;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_783_1;
    c_783_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxzz11x00zzz1xzxxz000x1xx11z10zxxxzzxxxzxzxxzxzxxxzzxxxzzxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

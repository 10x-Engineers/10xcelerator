class c_1033_1;
    integer i = -171;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1033_1;
    c_1033_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1x011zx11x1x10z1z1x0x100zx0zzx0zzxxzxzzzzxxzzzxzxzzxzxxxxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2715_1;
    integer i = -451;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2715_1;
    c_2715_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0xx1xz0xzzxx1100zxx0z0xzxx0xxxxzxzxzzxxzzzzzzxzzzxxxxxxzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

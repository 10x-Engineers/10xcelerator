class c_409_1;
    integer i = -67;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_409_1;
    c_409_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00xx111xx01xz1z10z11x1z111zxxzz0xxzzzzzzxzzzxxzxzzxzxzxxxzzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

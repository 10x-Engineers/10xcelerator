class c_2324_1;
    integer i = -386;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2324_1;
    c_2324_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1x0zxx1z11z1xxz111x1z1zzzxxz0zxxzxxxxxzxxzxzxzzzzzzxzzxxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2677_1;
    integer i = -445;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2677_1;
    c_2677_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xz11x1xxxxx1111z1x1z1xzz00zxx00xxzzzzzzxxxxxzxxzzzxzzzzxzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

package include_pkg;
  import uvm_pkg::*;
`include "uvm_macros.svh"



`include "Seq_item.sv"
`include "Relu_Sequence_item.sv"
`include "Seqr.sv"
`include "Sequence.sv"

`include "Driver.sv"
`include "Monitor.sv"
`include "Agent.sv"
`include "Passive_Monitor.sv"
`include "Passive_Agent.sv"

`include "environment.sv"
`include "Relu_Scoreboard.sv"
`include "Environment.sv"
`include "Conv_Scoreboard.sv"
`include "Test.sv"


endpackage
class c_1815_1;
    integer i = -301;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1815_1;
    c_1815_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zzzx1xz010x0110xxz100x0xz1011zzxxxzxzxzzxxxxzzxxxzzxzzxxzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_626_1;
    integer i = 626;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_626_1;
    c_626_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z0z0z0z0xzxx1z1xzz111z1xz0zzz0xzxzxxxzzzzxxzzzxzxzzzxzzxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_393_1;
    integer i = 393;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_393_1;
    c_393_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x111x010x0x110x1z0zz1z00xxx1zzzxzxzzzzxzxzxxxzzzxxxxxxxzzxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

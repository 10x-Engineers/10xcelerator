class c_2768_1;
    integer i = -460;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2768_1;
    c_2768_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zx010xx0x1z10xz01x111zxzz0110zxzxxxzzxxxxxzzzxxxxzzzxzxzzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

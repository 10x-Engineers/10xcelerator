class c_2498_1;
    integer i = -415;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2498_1;
    c_2498_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzxz10x01xxxxzzxz10z0z0z0zz1xz01xxxxxzzzzzxzxzxxxzxxzzxxzxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_703_1;
    integer i = 703;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_703_1;
    c_703_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z10x0xxzzzxx011z1zxzxx1zx0110z1xxxxzxxzxxxxxzxzxxzxzzxzzxxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_752_1;
    integer i = -124;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_752_1;
    c_752_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x1xx1zz1z1z000xzx001xxz1x0x1xzxzxxxxzzzxzzzxxzzzzxzzzxzxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

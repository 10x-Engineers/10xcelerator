class c_1570_1;
    integer i = -260;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1570_1;
    c_1570_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x110zzzxx110z1x0zz1x01xzxx0z0110xzzzzxzxxxzzzxzzzxxxxzzzzxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

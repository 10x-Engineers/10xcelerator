class c_1260_1;
    integer i = -208;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1260_1;
    c_1260_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0011x1zx0x01010zxxz1zxx000zz0z1xxzzxxxzzxzzxxzxxxzxzzxxxxxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

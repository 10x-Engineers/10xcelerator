class c_460_1;
    integer i = 460;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_460_1;
    c_460_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00100000zxzxxxx10001xz1zz1xx1x0zxxzzzxxxzxxxzzzxxxxxxzzxzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

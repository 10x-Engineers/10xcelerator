class c_1830_1;
    integer i = -303;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1830_1;
    c_1830_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxxx00x00zxx1xx1x10zz01xx0zx01zzzxxxxzzxzxxzxzxxxxxxxzxzzxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1077_1;
    integer i = -178;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1077_1;
    c_1077_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x10x1zxz0zz0x010z0111z11010x011xzzzzzzxxxxzxzzzxzxxzxxzxzzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1563_1;
    integer i = -259;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1563_1;
    c_1563_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1110x10z110xzz1z00xxxxx1xxzz0x1zzzxxxxxxxxxxxxxxzzzxzxzxxxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_128_1;
    integer i = -126;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_128_1;
    c_128_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x1z000z1z01zzx01zzxzxxxz1x010x1xxxxzzxxzzzxzxxxzzzxzxxzzzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

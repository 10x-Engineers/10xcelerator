class c_368_1;
    integer i = 368;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_368_1;
    c_368_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11000z0z01010xxz1x10xx0x1z0xxxxxxxxzzxzzxxzxxxxzxxzxzxxzzxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1187_1;
    integer i = -196;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1187_1;
    c_1187_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000xz11z0z1z110z010x00z10z0xzzxxzzzzxzzxxzxxxzzzzzxzxxzxxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

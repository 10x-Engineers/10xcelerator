class c_76_1;
    integer i = -74;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_76_1;
    c_76_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x101101z0xzx0zzzx0z00zz11zzzx1zxxzzxxzzxxzxxxzxzxzzzzxzzzxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_446_1;
    integer i = -73;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_446_1;
    c_446_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1z1z1x10z11111xz1xzzzxzz0z1zxxzzzzzxxxzxxzxzzzzzzxxxxxxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1136_1;
    integer i = -188;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1136_1;
    c_1136_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xzzx110xxzxz01z1xz10111x011z01zzxzzzzzzzxzxxxxzxzxzxxzxxzxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

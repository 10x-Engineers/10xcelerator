class c_476_1;
    integer i = -78;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_476_1;
    c_476_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z11zx01z1xz0zzxxzzxx0010x0x1zzzzzxxzxxxxzzzzxzxxzzzxzxxzxzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2429_1;
    integer i = -403;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2429_1;
    c_2429_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zz001xxz0z1x11z0xxz0xxzx011z11xzzzzzxxxzxxxxxxzzxzxxzzzzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

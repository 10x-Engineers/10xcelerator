class c_694_1;
    integer i = 694;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_694_1;
    c_694_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzz11xz0xz0x000xzzz1000xx01x01xxzzzzxxzxxzzzxxzxzxxxxzxxxxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1490_1;
    integer i = -247;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1490_1;
    c_1490_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010zz1x0x001z000x0x1010x01zzxxzxzxxzxzzxxzxzzxxzxzzzzxzzxzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

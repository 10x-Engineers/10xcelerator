class c_349_1;
    integer i = -347;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_349_1;
    c_349_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z111x011z011xz0z0zz111z1x0110z0xxxxzxxzxxxzxxzxzzxxzzzzzxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

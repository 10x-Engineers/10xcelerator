class c_958_1;
    integer i = -158;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_958_1;
    c_958_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1xz1z0x1111x11x1xzz111zxz0xx1zxxxzzzxxzxxzzxzxxzzxxxxxzxzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_868_1;
    integer i = -143;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_868_1;
    c_868_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z1x001x01011zzx1zx1000z1x11z10xzxxzxxzxxxxxzxxzxzzzxzzzzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

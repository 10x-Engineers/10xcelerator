class c_379_1;
    integer i = 379;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_379_1;
    c_379_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx10zz11zx110xzzz1z00z0x00zzz11zzxzzzzxzxxzzzzxzxzzzxxzzxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_429_1;
    integer i = -427;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_429_1;
    c_429_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx00zx01zz0z1zxz101xx01xzz10xz0xzxxxzxzxzxxzzxzzxzzzzxxxxzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

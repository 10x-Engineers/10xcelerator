class c_2750_1;
    integer i = -457;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2750_1;
    c_2750_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx1xzz000zz1z1zxxzx0z1zz01z1zx0xxzzxzxxzzxxzzzxxzzzzxxzzzzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

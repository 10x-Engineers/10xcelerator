class c_422_1;
    integer i = 422;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_422_1;
    c_422_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1x10010zzzx10110001x1x0111xx0zzxxzzzzxzzzzxzzzzxxzzzzxzzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

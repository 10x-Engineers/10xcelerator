class c_2937_1;
    integer i = -488;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2937_1;
    c_2937_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010011xx01001000111z0x110zx0z0z0zxzxzxzzxxxzzzxxxzzzzxzxzzxzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_953_1;
    integer i = -157;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_953_1;
    c_953_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0xx0x1xxx1x1xz0x1zx1xx00x1x010xzxxzzzzzzzzzzzxxzxxxxzxzxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

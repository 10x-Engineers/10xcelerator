class c_701_1;
    integer i = -699;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_701_1;
    c_701_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxz0xz10zz1x11001011x001x101xx1xzxxxxzzxzxxzzzzxzzxzzzzxxxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_429_1;
    integer i = -70;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_429_1;
    c_429_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx0x1z101zxx0x11x0z1z1zx00111zxxzxzxzxzzxxzzzxxzzxzxzzxzzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

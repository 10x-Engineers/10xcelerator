class c_2978_1;
    integer i = -495;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2978_1;
    c_2978_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00xx0xzxx110zzx111zx1zz11100x0xxzzzxxzxxzxxxxzxxzzzzzxzxxzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

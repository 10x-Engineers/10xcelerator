class c_1213_1;
    integer i = -201;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1213_1;
    c_1213_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zz1xz0zzzzz0xz1z00z10xxx01011zzxxxxxxzxzxxxzzxxxzxzzzxxxzzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_385_1;
    integer i = -383;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_385_1;
    c_385_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xx0zzxz10110z01xz1zx1z0x0xz0zx0zzzzxxzzxzxzzzzzxzxzzzxxzxzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2519_1;
    integer i = -418;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2519_1;
    c_2519_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010xxxxx01x100zx0z010xx000z10111zzxxzzxxzzzxxxxxxxzxxzzxxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

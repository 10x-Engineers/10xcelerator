class c_2038_1;
    integer i = -338;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2038_1;
    c_2038_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z1xzx1x11x0zxzzz1xx1zzx0x01x00zxxxxzxzzxxzzxxxxzxxzxzxzzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

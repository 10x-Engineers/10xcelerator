class c_403_1;
    integer i = 403;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_403_1;
    c_403_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11110z1zzzzxx10x00x0z000x0x01010xzzxxxxzxxzxzxxzxxzxzzzxxzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3362_1;
    integer i = -559;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3362_1;
    c_3362_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzz0xx110zxxxxx001zz10z01110zx0xxzzxxxxxzzzxzzzzzzzzzxxzzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_498_1;
    integer i = -81;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_498_1;
    c_498_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x011xx10xxxzxx0z1zzz1zx111xzz1xzxxxzzzxzxxxzzxzxxzxxzzzzxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2570_1;
    integer i = -427;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2570_1;
    c_2570_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1xz0xz0z011xz11z1z01z11x1zz111zxxzzxzzzxxxxxzzzxxxzxzzzxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

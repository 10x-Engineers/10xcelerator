class c_3282_1;
    integer i = -545;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3282_1;
    c_3282_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z0xz1x010x1x10zx010100x0zx0x10zzxxxxzzzxxzzzxzzxxxxzxzxxxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2954_1;
    integer i = -491;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2954_1;
    c_2954_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0x1xx0z1zxx1zxx1zxzxxzx01zzx0xzxxzxxxzxzxzzzxxxxzxxxzxzxzxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

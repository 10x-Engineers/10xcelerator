class c_1531_1;
    integer i = -254;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1531_1;
    c_1531_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzxx0zz001z0xxzz11x0z11xz111zx0zxxxxxxzxxzzzzzzxzxzxzzzzzxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3247_1;
    integer i = -540;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3247_1;
    c_3247_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xzz00z0xxx0zxzz11111x0xzzxz0zzzzxzzxxzzzxxxzzxzzxzxzzzzzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1353_1;
    integer i = -224;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1353_1;
    c_1353_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xxxz0x01xx10xz1z00zz0xx01xz1zxxzzxzxzzxxxxzxxxxzxxzzzzxxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

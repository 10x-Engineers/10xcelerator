class c_2966_1;
    integer i = -493;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2966_1;
    c_2966_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zxxx110z1111z000z11zx101x0zzz1xzzzxxzxxzzzzxzxzxzzzxxxzzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

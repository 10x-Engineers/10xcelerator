class c_544_1;
    integer i = 544;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_544_1;
    c_544_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz1z0100xzz110zx0111z1z1xxx01xxzxzzxxzzxzxzzxzzxxxzxzxxxzxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

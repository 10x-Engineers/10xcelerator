class c_626_1;
    integer i = -103;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_626_1;
    c_626_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxz010z0zxzxxx0x00zzzz1xxxxz10zxxzzzzxxzxzxxxxzxxzzxxzzxxxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_357_1;
    integer i = 357;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_357_1;
    c_357_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x111x10z1zzx01zxx1zxxz00z1000x1xzzxzzzxzxzxzxxxzzxzxzzzxxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

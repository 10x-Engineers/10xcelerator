class c_1204_1;
    integer i = -199;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1204_1;
    c_1204_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zx100z1010zxx0x01zxxzxz0xx001xxzzxzzzxxxzxzzxxxxxxzzxxxxzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_251_1;
    integer i = 251;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_251_1;
    c_251_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0100110zxxx000z0x11xx000xzzx0xzzzxxzzzzzzzzxzzzzzxzzxxxxzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2484_1;
    integer i = -412;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2484_1;
    c_2484_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xxzxz110xx11x0z0xz11zzz0xzzzx1xzxzzxxzzxzzzxzzzxzxxzxzxzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

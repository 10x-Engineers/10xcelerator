class c_805_1;
    integer i = -133;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_805_1;
    c_805_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xz000xxx1x1x1zzx1x010x1zxz0z10zxzzzxxxzzxxzzxzxxxzzzzxxxzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

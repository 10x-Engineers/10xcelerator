class c_788_1;
    integer i = -130;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_788_1;
    c_788_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x10xxxz000zxx00xzzzxzz11zxxxz0xxzzzzzzzxzxzzxzzxxzzxxxzxxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_628_1;
    integer i = -103;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_628_1;
    c_628_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xz000z11zzxzz0zzxzzzzxx10zx0xx0zzxzxxzzxxzzzzxzzxzzzxzxzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

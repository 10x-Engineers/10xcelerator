class c_2901_1;
    integer i = -482;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2901_1;
    c_2901_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzxx0zxzx1011000z0x0x1x1z001xz0xzzxzxzxzzxxxxzxxzxzxxxzxzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

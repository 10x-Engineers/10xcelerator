class c_818_1;
    integer i = -135;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_818_1;
    c_818_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zzzzx0x0xx0zzxx000zz1010zx1z11xxzxxzzzzzzzxzxzxxxzxzzzzxzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2942_1;
    integer i = -489;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2942_1;
    c_2942_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxz011zx0zx00z0111x1x1x1zz1z10zxzzzxxzxzxzzxxzzxxzzxzzzzxzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_134_1;
    integer i = -21;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_134_1;
    c_134_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0z1z1x0z1100z1x10zxxxxz0xx1xxxxzzzxxzxzzzxzxxzxzzzxxzzxxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

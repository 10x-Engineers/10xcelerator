class c_2101_1;
    integer i = -349;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2101_1;
    c_2101_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0x0zxxz1z0z0xzz10zzzz11xzxz011xzxxxxxzxxzzxxzxzxzxxzzzxzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3422_1;
    integer i = -569;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3422_1;
    c_3422_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z01z1z1101x1zz0zz1x11x0xzzzzz0xzxxxzxxxxzxzzxzzxxxxxxxxzxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

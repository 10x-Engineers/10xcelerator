class c_1566_1;
    integer i = -259;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1566_1;
    c_1566_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzz1x00zx1z0x0101x1x00z1zxzz10zzzxxxxxxzxxzzzzzxxxxxzxxxxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

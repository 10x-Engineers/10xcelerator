class c_1231_1;
    integer i = -204;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1231_1;
    c_1231_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zzz01z01zzx1zz1zx1x1xz0x0z1z01xzzxxxxxzxzzzzxxxxzzxxxxzzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

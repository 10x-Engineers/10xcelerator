class c_607_1;
    integer i = -100;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_607_1;
    c_607_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxz0x1xzxxxz000xzx101xx1101x10xzzxzxxzxxzzxzxxxxxzxzxxxzxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

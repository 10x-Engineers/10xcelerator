class c_3227_1;
    integer i = -536;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3227_1;
    c_3227_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xzx0z10xxzzzx0xx00z11zx10x100xxzxxzxxzxzxzzxzxzxxxzxzzzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1549_1;
    integer i = -257;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1549_1;
    c_1549_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1110z0x0xzz01x0110zz0xxzzx0zzxxzzxzzxxxxzzzxxzzzzzzzzxxxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_522_1;
    integer i = -520;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_522_1;
    c_522_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzz000010zzzxzx110xxxzz11z0zx00zxxxxxzxxxxxxzzzxzzxzxxxxxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2212_1;
    integer i = -367;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2212_1;
    c_2212_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx0x101zz0xz0z0zzx1x11z1xz010xxxxzzzzxzxxxzxxxxxxzzzzzzzxxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

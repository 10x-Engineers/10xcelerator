class c_418_1;
    integer i = 418;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_418_1;
    c_418_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1x0x0z1xz10zx10z0100z0z10110z0zxxxxzxzxxzxzzxxzzxzzzzxzxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3275_1;
    integer i = -544;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3275_1;
    c_3275_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0111zzxxxz0zxx1zzzzx0zxx11x01010xxxzxxzxzzxxxzzxzxxzzxzzzzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_851_1;
    integer i = -140;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_851_1;
    c_851_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzzx1z11xx11zz0zx1xzxx1x0x0zx00xzxzzzxxzzxzxzxxxzzxzxxxxzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_71_1;
    integer i = -10;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_71_1;
    c_71_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x011zz1zxxxzzx1xzx0001z011xxz1z1zzxxxzxzzzzzzxzzzzzxzzxzxzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

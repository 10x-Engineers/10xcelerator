class c_2612_1;
    integer i = -434;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2612_1;
    c_2612_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00z1xz11zz0zx1z10010zzz1z1z0100zxxxzzzxzzxzxxxzxxzxxzzzzxxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

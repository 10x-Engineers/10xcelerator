class c_181_1;
    integer i = -29;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_181_1;
    c_181_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0101xzzxzz11zz100xzz10zzzxzx1x1xzxzxzxxxzxxxxxzxxxzxxzzxzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1771_1;
    integer i = -294;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1771_1;
    c_1771_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10xz1zx011xz01xzz0zz1x0zx00xxzz1xzxxzzzzxzxxzzzzzxxzxzzzzzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

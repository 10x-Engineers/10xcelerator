class c_2784_1;
    integer i = -462;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2784_1;
    c_2784_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxx11111101x0xx11xz0x1zxz100xx10zxxxzzxzxzzzzzzxxzxzzxxzzzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

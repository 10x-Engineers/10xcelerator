class c_334_1;
    integer i = -54;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_334_1;
    c_334_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00000x011zxz101100xxzx1z01z01001zxzzxzzxzxzzxxxxxzzzzzzzxzxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

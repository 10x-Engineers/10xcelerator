class c_609_1;
    integer i = 609;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_609_1;
    c_609_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxxxx0xz1z110zx1z0z1xxx0zz00xx10xxzxzxxzzxzzzxzxzzzxxxxzzzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

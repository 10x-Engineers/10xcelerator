class c_142_1;
    integer i = 142;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_142_1;
    c_142_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00zxz0z1xxxxxxzxz01zz110100zzzzxzxxxzxxzzxzzzxzzxxxxxzzxzzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3210_1;
    integer i = -533;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3210_1;
    c_3210_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zx0xxxz111z000zz101xx010z11z10xzzxxxzxxzzzzzxzzzzzxzxxxzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_299_1;
    integer i = -48;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_299_1;
    c_299_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1001zzxz00z1z0zzxz0zxx0x011xzxxxzzxxxzxzxzzxxxzzzxzzxxxzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1781_1;
    integer i = -295;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1781_1;
    c_1781_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxxxxx11100x10xzzz101x01x01xx00zzxzzzxzzzzzzxzxzzxzzzzzxzzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

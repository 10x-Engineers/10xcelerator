class c_1003_1;
    integer i = -166;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1003_1;
    c_1003_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111xx1101x001zx01z1xxz0xxz0xxxzzzzxxxxxxxxxzzxxzxxxzzzxzzzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

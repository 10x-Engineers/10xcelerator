class c_2199_1;
    integer i = -365;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2199_1;
    c_2199_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x1zzz1zx00101zzzx101xz1xz1000x0zzxxxxxxxxxxxzzzxxzzzxxzzxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_338_1;
    integer i = -336;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_338_1;
    c_338_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xxz0x1z1x0xxzxxx001x0x0011z0zx0xxxxzzzxxxxzxzxxzxxzzxxzzzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_448_1;
    integer i = -446;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_448_1;
    c_448_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010x10x0110zz1z1111z0xx101111010xxzzzzxzzxxzzxzxzzxxzxxxxxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

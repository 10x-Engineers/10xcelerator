class c_3065_1;
    integer i = -509;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3065_1;
    c_3065_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzz110111z1z0x0z0z11x0x0xx0zz00zzxxzzxxzzzzxzxzxxzzzxzzxxzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

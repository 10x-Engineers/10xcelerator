class c_493_1;
    integer i = -491;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_493_1;
    c_493_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z1z1000011z1z1101zx10x0010zxz1zxxxzzzxxxzzxxxxxxxzxxxxzzxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

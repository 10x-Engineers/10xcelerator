class c_576_1;
    integer i = -94;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_576_1;
    c_576_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xx1z11000x1110z1z1x00zx1110x01zxxxxxxzxzxzxxzxzzxxzzxzzzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

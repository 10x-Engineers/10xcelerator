class c_506_1;
    integer i = 506;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_506_1;
    c_506_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx1xzx0xzxz010z0z11z0x1z1zx1zz0zzzxxzxzzzxzxzzzxzxxxzxzzxxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

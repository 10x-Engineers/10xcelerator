class c_20_1;
    integer i = -2;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_20_1;
    c_20_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzx1zzz011z0xx000z11xz00xzxzz11zzxxzxzxxxzxxzzxxxzzxxzzxxxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_520_1;
    integer i = -518;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_520_1;
    c_520_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1011z111z001xzzzzx11z0xzzxzxzzzxzxzxzxzxzzzxzzzzzzzxzxxxzzzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1361_1;
    integer i = -225;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1361_1;
    c_1361_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx01z00z10x0xxz0z0z0x1xzzx101zzzxxzzzzxzzxxxxzzxxzxzxxzxxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1643_1;
    integer i = -272;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1643_1;
    c_1643_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1xz010x00z1zx1xz00x00011x1x100xxxxxzzzzxxxxzxzxzxzzxxxzzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2892_1;
    integer i = -480;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2892_1;
    c_2892_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzx101x001z01z000000z0111zxx01zzzxzxxzzzxxzxxzxxxzzzxzxxzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1302_1;
    integer i = -215;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1302_1;
    c_1302_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x1zzx11xz01z0xzx1zx0z0xx11x0zzxzzzxzxzzxxxxzzzxxzzxzxxxzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

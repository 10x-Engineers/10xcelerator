class c_1718_1;
    integer i = -285;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1718_1;
    c_1718_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101zzx1z0z11011xz0z0xx011zx01111xxxzzzxzxxxxxzxzxxxxzxxzzzxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

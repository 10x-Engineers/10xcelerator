class c_744_1;
    integer i = -742;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_744_1;
    c_744_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx01xxz010zxzxxx011xxx110xzxx110zxzxzzxxzzzxzxzxzzxzzxxzzzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_287_1;
    integer i = -46;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_287_1;
    c_287_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z01z0xx00x1001x11xxx0zz1xzzxz0xzzxzxxxzxxzzxxxxxzzxxzzzzxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

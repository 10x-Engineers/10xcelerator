class c_2267_1;
    integer i = -376;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2267_1;
    c_2267_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x1zzz0zz0x000z1100zx01xz1x0z01zxzxxxzxxzzzzxxxzzzxzxzxzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

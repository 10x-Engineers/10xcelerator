class c_476_1;
    integer i = -474;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_476_1;
    c_476_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110x000z10zzx1zz1x0zz1z01x1x0z1xxxzzxzzxzxxxxzzzxxxzzxxxxxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2734_1;
    integer i = -454;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2734_1;
    c_2734_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0011zxzxzxxz0xz0zzx1xzx1zz1xzxzxxzzzxzzzxzxzxxzxzxzxxzzzzzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

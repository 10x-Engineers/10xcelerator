class c_1464_1;
    integer i = -242;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1464_1;
    c_1464_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xz01zzzzxz0z1z0zxxzx0z000x000zxxzzzzzxzxxxzzxxzxxxxzxzzxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

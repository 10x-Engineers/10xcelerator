class c_2249_1;
    integer i = -373;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2249_1;
    c_2249_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzz01zx00xxz0x0xz011x11011xxz11zxzzzzxxxzxxxxxxxxzzzxxxxxxzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1990_1;
    integer i = -330;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1990_1;
    c_1990_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz100zz1z0110xz1x1x11xz1zxx0xx1xzzzxzzxzzzxzxxzzxzzzzxxxzzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3017_1;
    integer i = -501;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3017_1;
    c_3017_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx101001z1xx0z00zzzz11zz0z1xz000zzzzxxxxzxxzzxxxzzzzxxxxxxxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

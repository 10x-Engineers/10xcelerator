class c_1224_1;
    integer i = -202;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1224_1;
    c_1224_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z001zz1xx1zx10xx1100xz0z1x10xxzzzzxxxzzzxxzzxzzxxzzxzxzzzxzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_525_1;
    integer i = -523;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_525_1;
    c_525_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10xzzxx0111z0xxxxzx1z0x0xz10x1xxxxxxxzxzzxxzzxxxxxxxxxxxzzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

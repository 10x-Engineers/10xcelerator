class c_2218_1;
    integer i = -368;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2218_1;
    c_2218_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00011x11xx1z10z01z0zz1zxzxx11110xxzzxzzxzxzxzzzzxzzzzzxzzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

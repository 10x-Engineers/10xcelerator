

interface small_if(input bit h_clk);


//int output_bits= 32; // fr time being hardcoding values 
//int input_bits =16;
        wire [32-1:0] output_port;
endinterface: small_if


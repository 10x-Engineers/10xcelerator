class c_2653_1;
    integer i = -441;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2653_1;
    c_2653_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xz0x0z01z011x1101zzx0xz0111x01xzzxzzzxzxxxzzxzzxzxzxzzxzxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_249_1;
    integer i = 249;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_249_1;
    c_249_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z001zx1xzz01010z1z10zz1zxzzzz0zzzzxzzzxxxzzzzxxxzzzxzxxxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_605_1;
    integer i = 605;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_605_1;
    c_605_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzx0xzz1xxx10z00z11zx1zxxzz0xz1xxzxzzxxzzxzxxzxxzxzzzxxxzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

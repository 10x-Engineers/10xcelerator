class c_1303_1;
    integer i = -216;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1303_1;
    c_1303_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111xzxx011z1101z1010x01010111000zzxxzzzzzxzxzzzzxzzzzzzxzzxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1347_1;
    integer i = -223;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1347_1;
    c_1347_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0zx0001z1001zz10000z0xzz1110x1xzzzzzxxzxzxxzzxxxzzxxxxxxxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

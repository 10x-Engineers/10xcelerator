class c_1046_1;
    integer i = -173;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1046_1;
    c_1046_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx010x1z01z001zz001111z0z1x0xz0zzzzxxzxzzxxxzxzxxzzzzzzzxxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_426_1;
    integer i = -424;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_426_1;
    c_426_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxxz11z1z0110xz110101011xz0x01zxxzxzzzxzxzxxxxxxzzzxxzxxzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

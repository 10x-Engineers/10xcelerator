class c_2449_1;
    integer i = -407;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2449_1;
    c_2449_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxxxz0z11xzzzz1x00z1zz111x1xz00zzzxzxxzxzzxzxxxxxxxzxzxxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_170_1;
    integer i = -168;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_170_1;
    c_170_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zz10xxz00x1zx10x01xxzz0x0z1z01xzzzzxxzxzzzxxzzzxxxzzzzzzzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_677_1;
    integer i = -675;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_677_1;
    c_677_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0zx1x0x011z1xzxxz100z11zxxzz1zxzxzzxzzzxxxzxzzzzxzxzxzzxzxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1897_1;
    integer i = -315;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1897_1;
    c_1897_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10z110111z0x1zzxzxzxxx0x1110z1zzzxzzzzzzzzzzxxzxzxzzxzzxxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_27_1;
    integer i = 27;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_27_1;
    c_27_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx011x0zxz1zxx0zzzx1x1xz01zxz111xzzxxxxxzxzzzzzxzxzxzzzxzzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_210_1;
    integer i = 210;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_210_1;
    c_210_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0x0101100110z0xx11z1z11xx0z101xxzzxxxzxxxzzzxzzzxxzzzzzzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

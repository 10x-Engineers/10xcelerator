class c_2117_1;
    integer i = -351;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2117_1;
    c_2117_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10110x00z00zxz01zzx0x1xxzxz10001zzzxzzxzzxzxxzxxxxxxxxzzzzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

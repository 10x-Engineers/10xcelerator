class c_502_1;
    integer i = -500;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_502_1;
    c_502_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxx001xx0xx0xx10z111zzxxzxx1xz0zzzxxzzzzxxxxxxxzxzxzzxzzxzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_741_1;
    integer i = -739;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_741_1;
    c_741_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xzzzxx0xxx1xz00000z101zz00zzx00xzxzzzzxzzzzzxzxxxzxxxzzxxzxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

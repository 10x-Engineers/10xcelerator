class c_278_1;
    integer i = -45;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_278_1;
    c_278_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzzx0101zx1z0z1z0z0zz0zz1z10zx01xzzzzzzxxxzzzzzxzxzzxxzxzxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

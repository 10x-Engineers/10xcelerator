class c_2115_1;
    integer i = -351;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2115_1;
    c_2115_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx101xzzxz010000zz000xzx0z111zzxzxxzxxxzxzxxzzxzxxzxxxxxxzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_395_1;
    integer i = -393;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_395_1;
    c_395_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0x10zzzx1x11xxx0100xx00x1100x1xxzxzzxxxxxxxxxzzxxxxzzxzzzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1685_1;
    integer i = -279;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1685_1;
    c_1685_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x01zx0x0101xx0z00x1z11x1zzz1xzzxzzxxzzxxzzzzzzxxzxzxzxxzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

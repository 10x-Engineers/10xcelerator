class c_2277_1;
    integer i = -378;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2277_1;
    c_2277_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10x011z1z0xxzx110zx0x00z0xz1000xzxzxxzxzxxzzxxxzzxxzzxxzzxzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_214_1;
    integer i = -34;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_214_1;
    c_214_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x1xx101z1zzxxx0zx1z1xx1x00x1xzzzzxxxxxzxxxzzzzxzxxzzzxzzxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

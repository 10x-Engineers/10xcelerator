class c_2895_1;
    integer i = -481;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2895_1;
    c_2895_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z000x11zxz1x1zz01zxzzzxxz0100xzzzzxxxzxzxxzzxzzxxzzxxzzzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_698_1;
    integer i = -696;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_698_1;
    c_698_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x110x01x111x11x0zxz1xzx110101zxzzxxzxxzxzxxxzzxxzxxxzxxzzxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1660_1;
    integer i = -275;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1660_1;
    c_1660_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "000z000z1z1zz0zzzxx11x1xx0xz0x0zxxzzxzxzzxzzxxxxzxxxxxzzxxzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

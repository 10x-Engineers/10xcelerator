class c_2818_1;
    integer i = -468;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2818_1;
    c_2818_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xz1zzxxz1x0100zx1z00xzxxz0zzx01zxzzzxzzxxxxxzzxxzzzzzzzzzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1818_1;
    integer i = -301;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1818_1;
    c_1818_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzx0zzx0z100z0x1xx0z1zx01zz0xz1zxzxzzxxzzxzxxxxxzzzxxxzzzzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2947_1;
    integer i = -490;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2947_1;
    c_2947_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x11zx1x101z01zxz11zx00zzzxxxz0zzxzxzzxxxzxzxzxxzxzxxxzxzxzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1126_1;
    integer i = -186;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1126_1;
    c_1126_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11x1xzxxxz011xxz00101x1x000zxxx0zzzzxxxzzxzzxxxxxxxzzzzxxzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3070_1;
    integer i = -510;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3070_1;
    c_3070_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xzxz0x00x1zxxxxx0x10011x0xxxz1xxzzzzzzxzzxxxxzxzzxxxxxzzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2490_1;
    integer i = -413;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2490_1;
    c_2490_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z11z1zxx11zz1z101xz1zx111xxxx0zzzxzzzzxxzxzzzxzzxxzxxxzzxzxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

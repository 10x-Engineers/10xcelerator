class c_2301_1;
    integer i = -382;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2301_1;
    c_2301_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx10z01011z10zxx11x101xx11zz01x0zzxzxzzxzxxzzzxzzzzxxzzxzxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

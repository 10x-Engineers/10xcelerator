class c_1515_1;
    integer i = -251;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1515_1;
    c_1515_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xxzxx0zx10xz00zx001xxx1111x0zzxzzzxxxzzxzxzxxzzxzzxzzzxzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_734_1;
    integer i = 734;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_734_1;
    c_734_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00xz00xxxz01x011xxxz111z0z00z0xzxzzxzxzxzxzxzzxxxxxzxxzxzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_507_1;
    integer i = 507;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_507_1;
    c_507_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1xx1xzx00zx10xzxx0xxxxx11zxx1zzzxzxzxzzxzxxzxxzzxzxzzxzxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1748_1;
    integer i = -290;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1748_1;
    c_1748_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz0x0100zz11x1zx0z0x0zz0010zz001xxxxzzzzzzzzzzxxzxzzzxxxzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

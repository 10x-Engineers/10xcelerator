class c_3381_1;
    integer i = -562;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3381_1;
    c_3381_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xx0xxxx1110x1zzzzxzxzx10xx0z01zzxzzxzxxzxxzzxxzxxxzxxzxzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

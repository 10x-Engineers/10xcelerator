class c_1405_1;
    integer i = -233;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1405_1;
    c_1405_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z0zxx0z10xzz0z10x1z0zxx1101x01xzxzzxzzxzzxxzzxzzxzzzxxzzxzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_422_1;
    integer i = -69;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_422_1;
    c_422_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xx1zxz1z0z1zzxz01110010xzzxxx0xzxxzxxxxxzzxxzxzzzzzzzzzxzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2967_1;
    integer i = -493;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2967_1;
    c_2967_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zx010xx001xxz0x1z1xz1zzzzx101zzxxzxxzzxxxzxzxzzzxxzxzzxxzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1892_1;
    integer i = -314;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1892_1;
    c_1892_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z00xzx1zx011x00x01101010zz110x1zzzxxzxzxxxzzzxxxxxzzzzxzxxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2675_1;
    integer i = -444;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2675_1;
    c_2675_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "011xz11x0z1xxzz11xzz0x0xz0z10101xxxzxxxzzxxzzzxxzxzzzzzzxxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_534_1;
    integer i = -532;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_534_1;
    c_534_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx1zzxxxx0zz0zxz1xzzxx1zx01x00z0xxzzxzxxxxzzzxxxxxxxzxzxxxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_333_1;
    integer i = -54;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_333_1;
    c_333_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001z101z1111x1zxzxxzx1x0zz00z0x0xzzxzxxzxzzzzzxzxxzxxzzxzxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_892_1;
    integer i = -147;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_892_1;
    c_892_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01z0x101xzz10zxzzzx0xzzz10xx0z10xzxzzxzxzxzzzxzxxxzzxzzzzzzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_33_1;
    integer i = -31;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_33_1;
    c_33_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx0xz1xzzz1110zxz1000x10zx1x00x1xzzzxzzxxxxxzxzxzxxxxzzxxxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1957_1;
    integer i = -325;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1957_1;
    c_1957_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xzx10x00x00x00111zx1z00000x1xxxzzzxxxxxxxzxxxzxzxzxzxzzxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

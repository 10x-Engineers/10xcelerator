class c_3125_1;
    integer i = -519;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3125_1;
    c_3125_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zzx1x10zx101100xxz0zxz001zzxz00xxxzzxxzxxxxzzxxxzxzzzzzxzzxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

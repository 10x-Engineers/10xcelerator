class c_189_1;
    integer i = -30;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_189_1;
    c_189_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "110z10111z11xx100x0xz0x011zz0x0zzxzzzxxxxxxzzzzxzzxxxzxxzxzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_662_1;
    integer i = -109;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_662_1;
    c_662_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z011xz0z10xxzx001x111z1zx0z1zzzxxzxzzzxzzzxzzzxzxxxzzzzzzzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

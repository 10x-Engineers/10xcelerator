class c_614_1;
    integer i = -101;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_614_1;
    c_614_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xz0x11xx100xzx111z10xxzz1xx1zxzzzzxzzzxxxxxzzxzxxzzzzxxxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1837_1;
    integer i = -305;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1837_1;
    c_1837_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11xzxx1zzzz11x0xx1001xxx1xxxzzz0xxxzzxxzzzxxxxzxxzxzzxxxxzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

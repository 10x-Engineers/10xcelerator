class c_2974_1;
    integer i = -494;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2974_1;
    c_2974_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z10xzzx0zzx1011x0z1zzxzxx1xz1000zzzzzxxzzzzzzzzzxxxzxzxzzzxzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2856_1;
    integer i = -474;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2856_1;
    c_2856_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzz1xxxz001z100xx01x0zzz1x001zz0zxzzxxxxzzxzxxxxzzxxxxzxxxxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1937_1;
    integer i = -321;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1937_1;
    c_1937_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1zxzxxxzz1xz0zz01xzz0x10x01zxxzzxxxxzxxzxzzxzzzzxxzzzzxzzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2508_1;
    integer i = -416;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2508_1;
    c_2508_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0x111xxx0xz1z010zz010x10x0zz0xxzzzxxzxzxzzzxxxzzzzzzxxzxxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

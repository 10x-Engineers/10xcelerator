class c_2158_1;
    integer i = -358;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2158_1;
    c_2158_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0001x00111x11xzz10x001xz1x10x1z0xxxzzzzxxxxxzxxxxzxxxxzxxxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

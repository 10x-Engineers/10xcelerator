class c_1439_1;
    integer i = -238;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1439_1;
    c_1439_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1100x001xz11x01z000010zx0zxz1zzxzzxxxzzxxzxxxzxzxzzzxxzxxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

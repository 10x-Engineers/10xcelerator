class c_483_1;
    integer i = -481;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_483_1;
    c_483_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xxzz1zzzxx0zx1011x11xzxz0z1z10zxxzxxxzzxxzzxxzxzxzzzxxzzxzxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3245_1;
    integer i = -539;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3245_1;
    c_3245_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z10xxzx0x1x1zxzxzxzxx1z1xxzxx1xxzzzzxxxzzzzzzzxzxxzxxzxxzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_366_1;
    integer i = -364;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_366_1;
    c_366_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x001xz110010zx0xz110xzxz1xz0zzzxxxzxzzxzzxxzxzxzxxxzxzzxxzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1722_1;
    integer i = -285;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1722_1;
    c_1722_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxxz101111zx1zx1x0z0z0xxx0xzz01xzzxzxxxxxzzxzzzzxzxxzzzxxxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_738_1;
    integer i = -736;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_738_1;
    c_738_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zz100011zxx10z1xzzz110zx1zz0zzxxzxzxzxzzxxxxxxxxxzxxxzxxxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2337_1;
    integer i = -388;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2337_1;
    c_2337_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z1zzxz1z1xx01xxz1zzzxz0x1zx0zzzzxxzxxxxxzzxzzzxxzxzxxxzxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

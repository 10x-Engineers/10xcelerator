class c_1108_1;
    integer i = -183;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1108_1;
    c_1108_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1z111x101xx0x10xzxx11111zxxz0xxzxxxxxxxxzxzzxzxzxzzxzzzxxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2125_1;
    integer i = -353;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2125_1;
    c_2125_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01x1xz01x1z101zx1001z0xxx1z0111xzzzxzxxxxxzxxzzxzzzzzzxzzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

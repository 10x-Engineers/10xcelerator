class c_3304_1;
    integer i = -549;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3304_1;
    c_3304_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0zx000z011xz0100z1z11zx00zxx0xxxxzxzzxzzzxxxxzxxxxxzzxzxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

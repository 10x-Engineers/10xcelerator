class c_731_1;
    integer i = 731;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_731_1;
    c_731_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00z1x0xz00zzz10xzzx101zxzzzx0z1xxzxzxzzzzzzxxxzxzxxxxxxzxxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

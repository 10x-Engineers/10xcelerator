class c_2650_1;
    integer i = -440;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2650_1;
    c_2650_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxzx011zz1100x1z11zxxz00x1xxx01zxzxxxzxzzxzxzxxzzzzxxzzzxxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2964_1;
    integer i = -492;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2964_1;
    c_2964_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "11zx11xzxzz1x1zx1xx0zz01zxzz0x01zxxzxxxxxxxzzxzxzxzxxzzzzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_764_1;
    integer i = -762;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_764_1;
    c_764_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zz00x11z1x111x11x10zz1z1zx111xxzzxxzzzxzxzzxzzxxxxzxzzzxxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1921_1;
    integer i = -319;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1921_1;
    c_1921_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xzx11xz01z10xzx1x01x1x1111z1zz0zxzxxxxxxzxxxzxxxzxzxxxxxxxxxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

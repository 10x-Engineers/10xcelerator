class c_1574_1;
    integer i = -261;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1574_1;
    c_1574_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z111101x0x0xzxzx0xx01zz0x1xxx0zzxxxxxzzzxzzzxzxzxxzxzxxxxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_754_1;
    integer i = -124;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_754_1;
    c_754_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxxz11xxx100101110z10xxzz00z11xxxxxzzxxzzzxxzzxxxxxzxxxzxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

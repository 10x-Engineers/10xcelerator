class c_1640_1;
    integer i = -272;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1640_1;
    c_1640_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x010zz11xzz10z11z11xx011zz011z0xzxzxxzzxzxzxxzzzzzzxzxzxxzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3097_1;
    integer i = -515;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3097_1;
    c_3097_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1x0zz1z110xz1z0zz0z0x0xzxzxx1zzzxxxzxxzxxxzxxxzxzxzzzzzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

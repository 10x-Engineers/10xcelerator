class c_1045_1;
    integer i = -173;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1045_1;
    c_1045_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01000001zz10z01x1101x10100z1011zxzxxzzxzzxzxxzxxzxxzxxzxzxxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_188_1;
    integer i = -186;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_188_1;
    c_188_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzx001z001zxz1zz1xx10z1xzz1z01xzxzzzzxzzzxxxzzxzxzzzzxzxzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

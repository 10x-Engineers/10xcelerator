class c_2771_1;
    integer i = -460;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2771_1;
    c_2771_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z001xxzz0z10z1zxxz100x1zxz01zzxxzxxxxzxzzzxzzzzxzzxxxxxzzzzzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

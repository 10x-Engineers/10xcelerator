class c_1900_1;
    integer i = -315;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1900_1;
    c_1900_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz010xzzz0111xzxz1x0111x1xz11zxzxxzzzzxzxxzxzxxxzxxzxzzxxxzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_274_1;
    integer i = 274;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_274_1;
    c_274_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zzzxxxx0x111xzxx1z0z11zx10z1zzzxzzxxzxxxxxzxxzzxzxzxxzxxzxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

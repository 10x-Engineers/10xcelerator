class c_24_1;
    integer i = 24;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_24_1;
    c_24_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxzxxx1x10z1x0zxz00010z0110x11xxzxzzzxzzxzxxzxzxxxxzxxzzzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3411_1;
    integer i = -567;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3411_1;
    c_3411_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1000z0zx1x10x111x0xzz10100z0100zxzzxzxxxzxzzzzzzxxzzxxxzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

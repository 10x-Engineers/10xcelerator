class c_932_1;
    integer i = -154;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_932_1;
    c_932_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx1z1z001xxxzzx0111xx1z11xx01zxxzzzzxzzzxxzzzzzzxzzzzxxzzxzzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

package include_pkg;
  import uvm_pkg::*;
`include "uvm_macros.svh"

`include "Sequence_item.sv"
`include "Seqr.sv"
`include "Sequence.sv"
`include "Driver.sv"
`include "Monitor.sv"
`include "Agent.sv"
`include "environment.sv"
`include "Environment.sv"
`include "Scoreboard.sv"
`include "Test.sv"
endpackage
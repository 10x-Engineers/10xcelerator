class c_1864_1;
    integer i = -309;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1864_1;
    c_1864_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x00zz00xxxx011zz0z1xxx1110x0xxzzzzzzzxxzzzzzxxzzzzxxzxzzzzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1170_1;
    integer i = -193;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1170_1;
    c_1170_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z100x11zx10z1xz0zx0x1101100x0110xxxxxzxxzzxxxxzzzzxxxxxzxxxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

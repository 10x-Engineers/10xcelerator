class c_1893_1;
    integer i = -314;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1893_1;
    c_1893_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx10zzxz0z001z01010z0z01xx1z00x0xzzzxzxxxxxzzxzxzzzxxzxxzxxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_348_1;
    integer i = 348;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_348_1;
    c_348_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1x1xzxx101x10xx11z0zx0011z01x1zzxzxxzxxxxxxzzxzxxxzzxxxzxzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_878_1;
    integer i = -145;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_878_1;
    c_878_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x10xzzxzzz1x1x0x010111x100001x0zzxxzxzzxzxxxzzzzzxzxxxxzxxxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2977_1;
    integer i = -495;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2977_1;
    c_2977_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101x1z10z0zxzzzzx01x110011zzzzxxzxxxzzzzzxzxxxxzzzxxxzzxzzxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

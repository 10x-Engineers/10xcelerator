class c_767_1;
    integer i = -126;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_767_1;
    c_767_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "001011z0z00z1x1001x1x0x1100x0z0zzxxzzxxxzzzzxxzzxzzzzzzzzxzzzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1399_1;
    integer i = -232;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1399_1;
    c_1399_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01xxxxz10zzz0zz00z00xx10x10xxxzxzzzzxzxzxxzxxzxzxxzzxzzxxxxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_841_1;
    integer i = -139;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_841_1;
    c_841_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x000011zxz111zxx0x10zx010z1z110zxxzzxzzxxxxxzxzzxzxzxzxxzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

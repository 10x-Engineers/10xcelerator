class c_39_1;
    integer i = -5;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_39_1;
    c_39_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00z0z0001z0xxz11010x0x1101x0110zxzxxzxzxxzxzxxxzxxzzzzzzxzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2731_1;
    integer i = -454;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2731_1;
    c_2731_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zx1z1z01zz01xz1xx01zx110zxz0xxxzzxxxxzzxzzzzzzzxxzzxxxxzzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_305_1;
    integer i = -49;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_305_1;
    c_305_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx1x010zx0zz0x0zxz11z1x00011xz0zzxxxxxxzxzzzzzzzzzzzzzzzzxzzxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

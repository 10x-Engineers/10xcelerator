class c_1085_1;
    integer i = -179;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1085_1;
    c_1085_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00zx0x00z10x0z0xx11xz0z1z1z0100zzxzxzxxzxzzzzxzxxxxxxzzxzzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2736_1;
    integer i = -454;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2736_1;
    c_2736_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00001z1x01zzz0x0x10x1z00010zxzzxzxxzxxzxzxxzxxzzxzzxxzxzxxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

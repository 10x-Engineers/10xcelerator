class c_51_1;
    integer i = 51;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_51_1;
    c_51_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1000zzzx11zxxzz0xzxzzz1xx01xxxxxxzzzzxzzxzzzxxxxxzzzxzxxzzxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1315_1;
    integer i = -218;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1315_1;
    c_1315_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz10z1100zx1x0zzzx10000zxz0x00z0zxzxzzxzzzzxzzzxzzxzxzzzxxxzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_625_1;
    integer i = -103;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_625_1;
    c_625_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xz0xz0xxzx1x1xz0z0010101000z10zzxxzxxxzzzzxxxzzxzxxxxzzxxxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_529_1;
    integer i = -87;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_529_1;
    c_529_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0z01xz1zxxxzx1xxz1z0z0xz011xxx1zzxzzxzzzxzzxzxxxzxxzxzzzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1044_1;
    integer i = -172;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1044_1;
    c_1044_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxzx101z001z0zxxzxzz1xxz1xx1zz1xzzxzxzxzzxxxzxxzxzzxzzxxzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1306_1;
    integer i = -216;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1306_1;
    c_1306_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz1111x0z0z0zx011100zxxzx11zx110zzxxxzxxxzzxzxzxxzzxzxxzxxzxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_554_1;
    integer i = -552;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_554_1;
    c_554_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1x010xx1xxz0zz0zxx00z0zz10x110zzzxzxxzzzzxzzxzxzzxxxxxxzxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1132_1;
    integer i = -187;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1132_1;
    c_1132_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxxzx110010xx10x0x001zxzz110xz1xzxxzzzzzxxxzzzxzxzxzxzxzzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2119_1;
    integer i = -352;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2119_1;
    c_2119_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "010z11zx0xxz110111x11zx0xx0xxxxxxzxxzxzxzxxxxxzxxxzzzzzzzxzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

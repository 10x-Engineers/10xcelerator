class c_250_1;
    integer i = -40;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_250_1;
    c_250_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxxx01x001xx1xx0z1xzx1zzxz1z00xxxxzxxxzzzxxxzzxzxzxzxxxxxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

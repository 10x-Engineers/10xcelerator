class c_1740_1;
    integer i = -288;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1740_1;
    c_1740_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z01x11zzz1zz10xxzzzz01z1xzzzz0x1zxxzxzzzzzxxzxxzxzxxxzzxxzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1536_1;
    integer i = -254;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1536_1;
    c_1536_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00xz0111xzzzzz011z01xxx1xzz0001zzzxxxzxxxxxzzzzzxxzzzxxxxxxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1899_1;
    integer i = -315;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1899_1;
    c_1899_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0zxz10z0xxx01zxzz0zzxz0x1x11x10xzxzxxzxxxzxzxxzzzxxzzzxzzzzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1269_1;
    integer i = -210;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1269_1;
    c_1269_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01z1x11z0100x000z1zz01z0110zxxzzzzxxzxzzzzxxzzzzxzzzzxxxzxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_39_1;
    integer i = -37;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_39_1;
    c_39_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z1z10z0xz111x1x0zzx1xxzxx0zxz1xxxzzzxxxzzzzxxzxzxzxzzxxxzzxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_628_1;
    integer i = 628;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_628_1;
    c_628_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zzzx111z01z0x0z10x01z10z00zzz0xxxxzxxzzzzzxzxxzxxzzzzzxxxxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

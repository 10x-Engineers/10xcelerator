class c_56_1;
    integer i = 56;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_56_1;
    c_56_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zx01xx01x010z0x0zzx0zzz100zxz1zzzxxzzxzxzzxzzzzxxxzzzzzzzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

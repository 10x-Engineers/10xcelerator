class c_588_1;
    integer i = -586;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_588_1;
    c_588_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x10x1zzzxx01100zz001x1z0xzzzx1zzzxxzzxzzzxxxzxzxxxzzzzxzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_775_1;
    integer i = 775;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_775_1;
    c_775_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10zzzz11x001x100zxz0xz01x0xzxxz1zzxxxxzxzzzxzxxzxxzzxzxzzxzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1338_1;
    integer i = -221;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1338_1;
    c_1338_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01xzx1zxxx0z0zx0x0x11x001x0xxxz1zxzzzzzxxzzxxxxxzxxzxzzxzzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1245_1;
    integer i = -206;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1245_1;
    c_1245_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x001z0z10x1x000xx101z0zxxzxxx1zxxxzxzzzzxzzzxzxzzzzzxzzzzxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2621_1;
    integer i = -435;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2621_1;
    c_2621_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z01xx011zzz1xx101z0001zx00000zzzxxzxxzzzxxxzxxzxzzzzxxzxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2005_1;
    integer i = -333;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2005_1;
    c_2005_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x001011000zx100010xz1zxzx1x1zxxxxxzzzzxzzxxzxxxxxxzxxzzxzzzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1542_1;
    integer i = -255;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1542_1;
    c_1542_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0z1zxzx1xx000z11xzzx100x10x101zzxzxzxzzzxzxxxzzzzxzzzxxzzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1351_1;
    integer i = -224;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1351_1;
    c_1351_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z0zzx11xz1z10x1110x011z00xxzx1zzxxzzzxxzxzzzxzxzxxxxzxzxzzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2382_1;
    integer i = -395;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2382_1;
    c_2382_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x011z1z10xx1xxxx01z0zxzzzxz0zzxxzxzxxzzxxzzxzzzxzxzxzzxzzxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3124_1;
    integer i = -519;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3124_1;
    c_3124_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xx111x0z1z0101x01x0zx00xx0xz10x0xzxzzxxxzzxzxxzxxzxxzzxxxxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

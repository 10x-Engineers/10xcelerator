class c_2820_1;
    integer i = -468;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2820_1;
    c_2820_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0zzz1z0zz1zx10zx1xzx11110110x1zxxxxxzzzxxzxxxxxzzxzzzxxxzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

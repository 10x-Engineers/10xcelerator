class c_3392_1;
    integer i = -564;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3392_1;
    c_3392_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zz011x0111z1z01x11z10zz1xz0zz001zxxxzzzxzzxxzzzxxxxzxzzxxxxzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_160_1;
    integer i = -158;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_160_1;
    c_160_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0zzxzzz10xz11z11zx0111x10x00x00zzxxzzxzzxxzzzxzxxzzzxzxxxzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

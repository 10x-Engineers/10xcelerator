class c_311_1;
    integer i = 311;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_311_1;
    c_311_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z111x001x1x00xzzzx00zzxx10xz0011zxxzzxxzxzxxxzzzxzxzxxzzxxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2483_1;
    integer i = -412;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2483_1;
    c_2483_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1zz100z0x10z01xx01x1x0xzz101z01xxxxzxzzzzzzxxxzzxxxxxzzxzxzxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_52_1;
    integer i = 52;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_52_1;
    c_52_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx100zzx00x0x01xxx1x1000zz10zz1zxxxxzzxxzzzxzxzzxzxzzzzzzxxxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_485_1;
    integer i = 485;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_485_1;
    c_485_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xzz1zzxzz1z0xz0zz011z01x0x100xzzxzxxxzzzzxzzzzzzxxxxxzzxxzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

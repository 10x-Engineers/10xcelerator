class c_812_1;
    integer i = -134;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_812_1;
    c_812_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x1x1xz100xz011z1x1z1xzx0x1z0zxx1zxxzzxzxzxxxzxxzzzzxxxxzzzzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_166_1;
    integer i = -164;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_166_1;
    c_166_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0x10x10xzz0xx1x011x110zz011zxz1xxzxxxxxzzxzxzzzxzxzzzzzzzxzxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

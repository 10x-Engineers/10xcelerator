class c_556_1;
    integer i = -91;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_556_1;
    c_556_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0xxx0x0xx0z11x100z1xz1x11101x1zzzzxzxxxxzxxzxzxxxzzxzzxxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_676_1;
    integer i = 676;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_676_1;
    c_676_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xz110zxxz0x1xxzx0x0zxxxzxx100xxzzzzzxxxxxxzzxzzzzxxxxzxzxxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1026_1;
    integer i = -169;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1026_1;
    c_1026_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z1x011xxx11100x1z100zxx0zz110z0zxzzxzzzxzxzxxxzxzzzzzxzxzxxxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

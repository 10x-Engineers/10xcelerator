class c_1226_1;
    integer i = -203;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1226_1;
    c_1226_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00x10xzx0100z111zzz10zzz011zxxx0xxzzzzzxxxzxxzzxxxzxxzzxzxxzzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_677_1;
    integer i = 677;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_677_1;
    c_677_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "101xz10x1xx1z100x1zxz1z10x000011zxxzzxxzxzzzxzzzxzxxzxxzzzxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_246_1;
    integer i = 246;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_246_1;
    c_246_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1zzxz001xzx0x11z0zz1zx00x1z100xzxzzxxzxzzzxzzzxxzzzxzxxzxzzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2091_1;
    integer i = -347;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2091_1;
    c_2091_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x11xxxx0xx1xx1x00100x11zz111zzzxxxxzxxzzxxxxzxxxzzzxxzxzxzzxzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_220_1;
    integer i = -35;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_220_1;
    c_220_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z111zx010z1xz0x1xzz0010z010xx1z0xzzzxxzxxxxzxzzzzxzxzxzxzxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

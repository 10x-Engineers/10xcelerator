class c_1469_1;
    integer i = -243;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1469_1;
    c_1469_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0z0xxz00zzzx0xz1z0xx11zxz00100x1zxxxxxxxzzxzzxxzzxxzzxxxzxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_290_1;
    integer i = 290;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_290_1;
    c_290_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xzzxx10x0z01001zz0111z1xx1010zxzxzxxzxxxxzzzzxxxxzxzzxzxzxzzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_3085_1;
    integer i = -513;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3085_1;
    c_3085_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1x0x001z1xx10x1z01101x1z0xzz0xzxxzxxxzxxzxzxzzxzxxxzzzzxxxxxzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

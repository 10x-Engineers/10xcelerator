class c_1055_1;
    integer i = -174;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1055_1;
    c_1055_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "111zzzx01x1x0zzzxzz0zzz11x1zzzxzxxxzzxzzzzzzxzzzzzxzzxzzzxzxzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_666_1;
    integer i = -109;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_666_1;
    c_666_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z1zzz10z1zzxxxz100x1x110xx0x11zxzxzzxzzxxxzzzzzzxzxxzzxzzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_653_1;
    integer i = 653;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_653_1;
    c_653_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00xzz0xx011z010x1z1x000xxz0zzzx0zzxzzzxxzzzzzxzzzxzxzzxzxxxzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_595_1;
    integer i = -98;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_595_1;
    c_595_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "01x10zz10zxzzz0xxx0xxxxx1x11100zzzzzxxxzzxxzxzxxxxxxzxxzxxzzzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

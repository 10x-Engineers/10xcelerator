class c_1664_1;
    integer i = -276;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1664_1;
    c_1664_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "0xxzz110zzx0z0x1x0zxx01xxzxzzz10zxzzzxzzxxxzzxzxzzxzxxxxxxzzxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

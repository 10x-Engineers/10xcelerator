class c_245_1;
    integer i = -243;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_245_1;
    c_245_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "xz1zxxz1xzz1xzx0xz1xx0xx11zz00x0xxzzxxzzzzxzxzzxxzzzxzxxxxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_872_1;
    integer i = -144;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_872_1;
    c_872_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xx011x11001x011011xz001x011z00zxzxzzxzxzxxzzxxxzzxxzzxxxzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

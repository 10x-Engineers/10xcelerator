class c_391_1;
    integer i = 391;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_391_1;
    c_391_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1001xz00xxxz1x1x1xzz110x1xzxzzxxxzxxxxzxxxxzxxxxxzzzzxxzzxzxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_543_1;
    integer i = -541;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_543_1;
    c_543_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00x0x0xx0xxz101011xx101z0z01z0zzxzxzzzzzxxxxxxzzxxxxzxzzzzxxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

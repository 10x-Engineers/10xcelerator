class c_676_1;
    integer i = -111;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_676_1;
    c_676_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zzx010z01x10x01x0x11zzzxxx101xxzzzzxzxzxxzzzzxzxxxxxzzzxxxxzxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_14_1;
    integer i = -1;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_14_1;
    c_14_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1xzz1xx1x0xz0x1101x0zxz1zzx1x01xzxzxzxxxxxzzxzzzxzzxzxxzxxzxxxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

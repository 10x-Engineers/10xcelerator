class c_2160_1;
    integer i = -358;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2160_1;
    c_2160_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z110x1xx0zxxxz11100xx0zz10xzz0x0zzxxxxxzxxzxxzzzxzxzxzxzxxxxzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

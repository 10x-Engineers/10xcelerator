class c_342_1;
    integer i = -340;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_342_1;
    c_342_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z00zzzzx1101xxzx1x0xx00xz0xz0100zzxzxzxxzxzxzzxzzxzzzxzxzzxzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

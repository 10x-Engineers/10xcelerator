class c_2376_1;
    integer i = -394;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2376_1;
    c_2376_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zxzxz1x0x00000zz101xx01xzxz1xx10zxzxzxxzxzxxzxzzxxxxzzxxxzzzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

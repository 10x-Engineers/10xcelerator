class c_1661_1;
    integer i = -275;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1661_1;
    c_1661_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x10x01110x00z00x101xz01zxzz11x1zzzxzzzxxzxxxxxxxzxxxxxxzxzxxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_486_1;
    integer i = -484;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_486_1;
    c_486_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "00z0xx00x10zxxx11x00z10000xzzxz0xzzzxxzxzzzxzzxzzxzzxxzzzzzxxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

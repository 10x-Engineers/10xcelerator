class c_216_1;
    integer i = -34;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_216_1;
    c_216_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z1x0zxx1z0xzzx01z00011xz01zxx1zxzzxzxxxxxxxzxxxzxzxzzzzzxxxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_578_1;
    integer i = -576;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_input_port == i);
    }
endclass

program p_578_1;
    c_578_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "10z1z01xz1zx1zxxx0zzx0xz1xzxzzx1xxzxxzxzxxzxxzzxzxxzzzzzxzzzzzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

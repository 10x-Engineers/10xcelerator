class c_3321_1;
    integer i = -552;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_3321_1;
    c_3321_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z0z00z10z11xxx011xxxzz1xz10x101zzxzzxzxzxxxxxzxxzxzxxxxxzxzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_1348_1;
    integer i = -223;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_1348_1;
    c_1348_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zx01zxzz00x000z0z0001x10xz1z00zzzzxxzzxzzxxzxxzzzxxxxxxxzzzxzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2611_1;
    integer i = -434;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2611_1;
    c_2611_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx1x00z100z1xz01100xz1x0xx10xz1zzxxxxzzxzzzxzzzzxzzxxxxzzxxxzxxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_732_1;
    integer i = 732;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_732_1;
    c_732_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzxx1xz0zz1z0010zz0xz10zz00x00zxxxxxzxxzxzxxxzzxzzxzxxxxxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_162_1;
    integer i = 162;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_162_1;
    c_162_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1z11111xz0x1101x110zzz00x1x101z1xzxxxxzxzzzxxzxzzxzzxzzxxzxxzzzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_675_1;
    integer i = -111;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_675_1;
    c_675_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xzxx101x0zxxzx1zx011zzxx01xzz1xzxxxxxzxzxzzzxxxxzxxxxzzxxzzxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_2246_1;
    integer i = -373;
    rand bit[15:0] tr_Input_Pixel; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       (tr_Input_Pixel == i);
    }
endclass

program p_2246_1;
    c_2246_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x01z1z011xx10xx110x0x1z1xxzz0010zxzxxxzzxzxxxzzxxzxxxzxzxzxxxzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram

class c_429_1;
    integer i = 429;
    rand bit[15:0] tr_input_port; // rand_mode = ON 

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (sequence.sv:17)
    {
       ((tr_input_port[15:13]) == i);
    }
endclass

program p_429_1;
    c_429_1 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z0xzxx00z1x0x01111xz0z1zzzxzz1xzzzxzzzxxxzzzzzzzxxzzzxxxzzxzxzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
